��]      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�_sklearn_version��1.5.1�ub�n_estimators�Kd�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK*�verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hNhG        �feature_names_in_��joblib.numpy_pickle��NumpyArrayWrapper���)��}�(�subclass��numpy��ndarray����shape�K���order��C��dtype�h-�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�
allow_mmap���numpy_array_alignment_bytes�Kub�cnumpy.core.multiarray
_reconstruct
q cnumpy
ndarray
qK �qc_codecs
encode
qX   bqX   latin1q�qRq�qRq	(KK�q
cnumpy
dtype
qX   O8q���qRq(KX   |qNNNJ����J����K?tqb�]q(X   PclassqX   SexqX   AgeqX   SibSpqX   ParchqX   FareqX   Embarkedqetqb.��       �n_features_in_�K�
_n_samples�M��
n_outputs_�K�classes_�h))��}�(h,h/h0K��h2h3h4h6�i8�����R�(K�<�NNNJ����J����K t�bh<�h=Kub�����               ��       �
n_classes_�K�_n_samples_bootstrap�M��
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJf��_hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4h6�f8�����R�(KhHNNNJ����J����K t�bh<�h=Kub��������������              �?��       hJ�numpy.core.multiarray��scalar���hGC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub���       �k      K��R�}�(hK�
node_count�M9�nodes�h))��}�(h,h/h0M9��h2h3h4h6�V64�����R�(Kh:N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(hqh6�i8�����R�(KhHNNNJ����J����K t�bK ��hrh}K��hsh}K��hthVK��huhVK ��hvh}K(��hwhVK0��hxh6�u1�����R�(Kh:NNNJ����J����K t�bK8��uK@KKt�bh<�h=Kub���       d                    �?���*1�?�           8�@               -                 �|Y=@���	���?^            �b@                                   �?��0u���?*             N@                                  �2@@4և���?             <@                                   �?r�q��?	             (@                               pFt*@"pc�
�?             &@        ������������������������       �                     @                                   �?�q�q�?             @       	       
                      @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@                                   @     ��?             @@        ������������������������       �                      @               &                    �?      �?             >@                                    @b�2�tk�?             2@                                �U�X@      �?              @                                �}S@r�q��?             @        ������������������������       �                     @                                  �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @               !                 ��Y&@���Q��?             $@                                ���@z�G�z�?             @        ������������������������       �                     �?                                   @@      �?             @                                 �5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        "       %                    �?���Q��?             @        #       $                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        '       ,                   �7@�q�q�?             (@       (       )                    �?�q�q�?             @        ������������������������       �                     @        *       +                 ��&@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        .       U                    �?��9܂�?4            @V@       /       P                    �?rr�J��?)            �R@       0       E                     �?V��z4�?"             O@       1       D                    P@�eP*L��?            �@@       2       5                    �?���>4��?             <@        3       4                 �iE@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        6       A                    C@     ��?
             0@       7       8                 ��";@�θ�?             *@        ������������������������       �                     �?        9       @                 @�Cq@r�q��?             (@       :       ?                 �|�=@�C��2(�?             &@       ;       >                 ��2>@z�G�z�?             @        <       =                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        B       C                 ��Y>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        F       O                 �|�=@\-��p�?             =@       G       H                    �?����X�?             ,@        ������������������������       �                      @        I       J                     @r�q��?             (@        ������������������������       �                      @        K       L                 ���@z�G�z�?             $@        ������������������������       �                      @        M       N                   @@      �?              @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     .@        Q       T                    �?r�q��?             (@       R       S                   �H@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        V       _                    �?�q�q�?             .@       W       X                   @D@      �?              @        ������������������������       �                      @        Y       ^                   @N@�q�q�?             @       Z       ]                      @      �?             @       [       \                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        `       a                     �?؇���X�?             @       ������������������������       �                     @        b       c                    :@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        e       2                   @��J���?f           ��@       f       y                   �0@n��6g�?V           ��@        g       n                     @�������?             F@       h       i                    �?HP�s��?             9@       ������������������������       �        
             *@        j       m                     �?r�q��?             (@        k       l                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        o       x                     @p�ݯ��?             3@       p       q                    /@      �?             0@       ������������������������       �                     "@        r       w                 pFD!@և���X�?             @       s       t                    �?      �?             @        ������������������������       �                     �?        u       v                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        z       �                 ���'@J��8�M�?8            @       {       |                 ���@�����?�            �o@        ������������������������       �                     >@        }       �                    �?�-��}x�?�            �k@        ~       �                    �?�Ƀ aA�?#            �M@              �                    �?�`���?            �H@        �       �                    �?z�G�z�?
             .@       �       �                 �|�9@$�q-�?	             *@        ������������������������       �                     �?        �       �                  ��@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        �       �                    3@ҳ�wY;�?             A@        �       �                    �?r�q��?             @       �       �                   �1@z�G�z�?             @        ������������������������       �                     �?        �       �                 ��!@      �?             @       �       �                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                     @      �?             <@        �       �                   �J@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                   �9@�}�+r��?
             3@        ������������������������       �                     $@        �       �                 @3�@�����H�?             "@       �       �                 �?�@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?ףp=
�?             $@       �       �                 P�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?ĴF���?f            �d@       �       �                   �>@�-���?`            `c@       �       �                 ���@�5̾�?O            �_@        ������������������������       �                     �?        �       �                 @3�@|�(��?N            �_@       �       �                   �<@�n���?+             R@       ������������������������       �                    �A@        �       �                 �|Y=@$G$n��?            �B@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��@�FVQ&�?            �@@       ������������������������       �                     8@        �       �                 �Y5@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                     @PN��T'�?#             K@        �       �                    5@�C��2(�?             &@       �       �                   �2@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 pf� @�T|n�q�?            �E@        �       �                 ��) @���y4F�?             3@       �       �                   �4@r�q��?             2@        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     ,@        ������������������������       �                     �?        �       �                 ���"@      �?             8@        �       �                    9@$�q-�?             *@       ������������������������       �                     $@        �       �                 �|Y<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �<@"pc�
�?             &@       ������������������������       �                      @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     <@        ������������������������       �                     "@        �                        x#J@L����?�            `n@       �       �                    �?�+Fi��?{             g@        �       �                 03�;@�M;q��?1            �R@       �       �                    �?�z�6�?(             O@        ������������������������       �                     @        �       �                   �2@x��}�?$            �K@        �       �                     @և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?     ��?              H@        �       �                   �+@���7�?             6@        �       �                    �?ףp=
�?             $@       �       �                    B@�����H�?             "@       ������������������������       �                     @        �       �                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             (@        �       �                    �?�	j*D�?             :@       �       �                    D@�ՙ/�?             5@       �       �                    �?�q�q�?             2@       �       �                 �|Y>@ףp=
�?             $@       ������������������������       �                     @        �       �                   �@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 0339@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                   @F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @�	j*D�?	             *@        ������������������������       �                     @        ������������������������       �                     "@        �                           �?�aV����?J            @[@        �       �                 �|�<@�X���?             F@        ������������������������       �                     @        �                         �>@��Sݭg�?            �C@       �                         �J@�G��l��?             5@       �                         `G@j���� �?
             1@       �                         @=@��S���?             .@       �       �                 03:@�q�q�?             (@        ������������������������       �                      @        �       �                 03k:@      �?             $@        ������������������������       �                     @        �                         �C@����X�?             @        �                        �|�?@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             2@                                 �?���Ls�?0            @P@                                �?��GEI_�?.            �N@       	      
                �|=@(N:!���?            �A@        ������������������������       �        
             1@                                 �?�<ݚ�?             2@                               �*@������?             1@                               �F@�	j*D�?             *@                             �|�=@X�<ݚ�?             "@        ������������������������       �                     �?                                 @@      �?              @        ������������������������       �                     �?                                �C@և���X�?             @                               �A@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     :@                                 �?      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 �?�e�,��?             �M@       ������������������������       �                     =@               1                   �?d��0u��?             >@       !      ,                    @J�8���?             =@       "      #                `�iJ@�z�G��?             4@        ������������������������       �                      @        $      +                  �D@�<ݚ�?
             2@       %      &                   �?���|���?             &@        ������������������������       �                     @        '      *                  �B@�q�q�?             @       (      )                   A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        -      0                �|�>@X�<ݚ�?             "@       .      /                �|�;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        3      8                   @���7�?             6@        4      7                   �?�����H�?             "@        5      6                   @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             *@        �1       �values�h))��}�(h,h/h0M9KK��h2h3h4hVh<�h=Kub�����`l����??'��d�?�m�PM��?ɟWY��?""""""�?�������?�$I�$I�?n۶m۶�?UUUUUU�?�������?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?�������?333333�?              �?      �?                      �?              �?              �?      �?      �?              �?      �?      �?9��8���?�8��8��?      �?      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?333333�?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?         ��G?��?�.p��?Z7�"�u�?L�Ϻ��?2�c�1�?�s�9��?t�E]t�?]t�E�?n۶m۶�?I�$I�$�?UUUUUU�?�������?      �?                      �?      �?      �?ى�؉��?�؉�؉�?              �?�������?UUUUUU�?]t�E�?F]t�E�?�������?�������?      �?      �?      �?                      �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        a����?�{a���?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        �������?�������?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        UUUUUU�?�������?F]t�E�?]t�E�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        _Xw
=�?CO���?�M1j���?�d�+H�?/�袋.�?t�E]t�?{�G�z�?q=
ףp�?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?Cy�5��?^Cy�5�?      �?      �?              �?�$I�$I�?۶m۶m�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        !�B!�?���{��?TqК3�?�:��1��?      �?        ;Ӹ�Qg�?���b�?~ylE�p�?'u_�?����S�?և���X�?�������?�������?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?UUUUUU�?�������?�������?�������?              �?      �?      �?      �?      �?              �?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        �5��P�?(�����?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?�������?�������?              �?      �?              �?        E�JԮD�?ە�]�ڵ?=���?�qa�?����x�?���p8�?              �?-˲,˲�?��i��i�?r�q��?r�qǱ?      �?        к����?���L�?      �?      �?              �?      �?        >����?|���?      �?        9��8���?�q�q�?              �?      �?        &���^B�?h/�����?]t�E�?F]t�E�?�������?�������?      �?              �?      �?      �?        ���)k��?6eMYS��?6��P^C�?(������?�������?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?        /�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        #e�����?�5?,R�?���,d!�?����7��?ƒ_,���?�6�i��?�Zk����?J)��RJ�?              �?A��)A�?pX���o�?�$I�$I�?۶m۶m�?              �?      �?              �?      �?F]t�E�?�.�袋�?�������?�������?�q�q�?�q�q�?              �?      �?      �?      �?                      �?              �?              �?;�;��?vb'vb'�?�a�a�?�<��<��?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?vb'vb'�?;�;��?              �?      �?        \������?������?]t�E�?�E]t��?              �?�|˷|��?�i�i�?1�0��?��y��y�?ZZZZZZ�?�������?�������?�?�������?�������?      �?              �?      �?              �?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?                      �?              �?      �?              �?        �����?z�z��?�d����?;ڼOqɰ?|�W|�W�?�A�A�?      �?        9��8���?�q�q�?xxxxxx�?�?vb'vb'�?;�;��?r�q��?�q�q�?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?              �?              �?              �?              �?      �?              �?      �?        _[4��?�pR���?              �?DDDDDD�?wwwwww�?�rO#,��?|a���?ffffff�?333333�?              �?9��8���?�q�q�?]t�E]�?F]t�E�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        r�q��?�q�q�?�������?UUUUUU�?              �?      �?                      �?              �?�.�袋�?F]t�E�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�=�KhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       j                    �?\AK"���?�           8�@               e                 ���Q@d��4a�?�             n@              ^                    @r��p���?z            �h@                               `f�$@Zb��'��?o            `f@                                   3@�Q����?             D@        ������������������������       �                      @                                 ��@�s��:��?             C@              	                    8@8����?             7@        ������������������������       �                     @        
                        ���@j���� �?             1@        ������������������������       �                     @                                  �9@�θ�?             *@        ������������������������       �                     �?                                ���@r�q��?
             (@        ������������������������       �                      @                                   �?z�G�z�?             $@                               �&B@      �?              @                                  �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                �Y5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                �|Y>@��S�ۿ?	             .@       ������������������������       �                     *@                                 SE"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               S                   �E@�S^�,�?T            `a@              H                 039@"pc�
�?J            @^@               1                    �?��M���?+             Q@        !       0                    �?���|���?             6@       "       '                    �?X�<ݚ�?             2@        #       $                     @      �?              @        ������������������������       �                     @        %       &                 03�-@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        (       /                 �|�<@      �?             $@       )       .                   �-@      �?              @        *       -                    �?���Q��?             @       +       ,                 �&�)@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        2       ;                    �?�5��
J�?             G@       3       8                   @B@ܷ��?��?             =@       4       5                     @$�q-�?             :@       ������������������������       �                     2@        6       7                 ��&@      �?              @        ������������������������       �                      @        ������������������������       �                     @        9       :                   �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        <       =                     @��.k���?
             1@        ������������������������       �                      @        >       ?                    �?���Q��?	             .@        ������������������������       �                     �?        @       G                 ���1@և���X�?             ,@       A       D                    �?z�G�z�?             $@        B       C                 �|�;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        E       F                    0@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        I       N                    �? �h�7W�?            �J@       J       K                     @@�E�x�?            �H@       ������������������������       �                    �G@        L       M                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        O       P                    @      �?             @        ������������������������       �                     �?        Q       R                   �6@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        T       ]                    �?b�2�tk�?
             2@       U       V                   �G@���|���?             &@        ������������������������       �                      @        W       \                    �?�<ݚ�?             "@       X       [                     �?�q�q�?             @       Y       Z                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        _       `                    @�<ݚ�?             2@        ������������������������       �                     @        a       b                 ���3@�q�q�?             (@        ������������������������       �                     @        c       d                    @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        f       g                  "�b@���7�?             F@       ������������������������       �                     @@        h       i                    !@r�q��?	             (@        ������������������������       �                      @        ������������������������       �                     $@        k       l                    �?�ְ�Hj�?)           `}@        ������������������������       �                     @        m       �                     �?l����~�?$           �|@        n       u                   �;@Ȩ�I��?A            �Z@        o       t                  "&d@      �?             0@       p       s                    �?����X�?
             ,@       q       r                   �8@�q�q�?	             (@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        v       �                    �?z�G�z�?5            �V@       w       �                    �?b�h�d.�?*            �Q@        x       �                   �F@z�G�z�?             4@       y       �                 p�w@�q�q�?	             (@       z       �                   @C@z�G�z�?             $@       {       �                 ��2>@�����H�?             "@        |                           �?z�G�z�?             @       }       ~                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �>@�J�4�?             I@       �       �                   �<@r֛w���?             ?@        ������������������������       �                     �?        �       �                 ��$:@�������?             >@        ������������������������       �                     $@        �       �                 X�,@@��Q��?
             4@        ������������������������       �                     @        �       �                 03k:@��S���?             .@        ������������������������       �                      @        �       �                 `f�<@�n_Y�K�?             *@       �       �                   �K@�q�q�?             (@        �       �                    H@      �?              @       ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     3@        �       �                    �?�z�G��?             4@       �       �                   @G@և���X�?             ,@       �       �                 `f�N@���!pc�?             &@       �       �                  x#J@      �?             @        ������������������������       �                      @        �       �                 `�iJ@      �?             @        ������������������������       �                      @        �       �                    A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �                         @@@�D�d@6�?�            Pv@       �       �                 ��K.@Pe6�p�?�            �p@       �       �                    ,@���d���?�            `i@        ������������������������       �                      @        �       �                    �?t�e�í�?�             i@        �       �                     @ȵHPS!�?             :@        ������������������������       �                      @        �       �                 ��� @      �?             8@       �       �                 �|Y=@؇���X�?             5@        �       �                    �?և���X�?             @       �       �                    ;@      �?             @       �       �                 ��y@���Q��?             @        ������������������������       �                     �?        �       �                   �6@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     @        �       �                 �|�=@4����Y�?t            �e@       �       �                    �?�G�z.�?i             d@       �       �                   �<@ �h�7W�?h            �c@       �       �                    �? �q�q�??             X@       �       �                 0S5 @XB���?9            �U@       �       �                 @3�@�X�<ݺ?#             K@       �       �                    �?@�E�x�?            �H@        ������������������������       �                      @        �       �                   �7@`Ql�R�?            �G@       ������������������������       �                     ?@        �       �                 ���@      �?             0@        �       �                   �8@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             (@        �       �                    3@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �@@        �       �                   �4@�����H�?             "@        �       �                    3@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���@�[|x��?)            �O@        ������������������������       �                     2@        �       �                     @�����H�?            �F@        ������������������������       �                      @        �       �                  sW@X�EQ]N�?            �E@        �       �                 ��@�<ݚ�?
             2@       �       �                 �|Y=@؇���X�?             ,@        ������������������������       �                     �?        ������������������������       �$�q-�?             *@        ������������������������       �      �?             @        �       �                 �|Y=@`2U0*��?             9@        ������������������������       �                     �?        �       �                 ��) @ �q�q�?             8@       ������������������������       �                     4@        �       �                 pf� @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                     @z�G�z�?             .@        ������������������������       �                     @        �       �                   �>@�q�q�?             "@        �       �                 �̌!@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��.@�̚��?"            �N@        ������������������������       �                     @        �                          �?P̏����?!            �L@       �       �                    �?�q�q�?             H@        �       �                     @�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        �                           �?���@��?            �B@       �       �                    �?      �?             8@        �       �                    �?�eP*L��?             &@        ������������������������       �                     �?        �       �                 �T�C@      �?             $@        ������������������������       �                     @        �       �                    ;@r�q��?             @        ������������������������       �                     @        �       �                    >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     @$�q-�?             *@        ������������������������       �                     @        �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?                                 @8�Z$���?	             *@                                 @�q�q�?             @                                 @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        	      
                  �D@�L��ȕ?6            @W@       ������������������������       �        !            �M@                                @E@г�wY;�?             A@                                  @z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     =@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������T1�m��?X�]$���?�֖�֖�?�������?e
�d�?��3�M��?��¨N�?x����X�?�������?ffffff�?              �?��k(��?�k(���?8��Moz�?d!Y�B�?              �?ZZZZZZ�?�������?      �?        �؉�؉�?ى�؉��?      �?        UUUUUU�?�������?              �?�������?�������?      �?      �?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?      �?      �?                      �?�������?�?      �?              �?      �?              �?      �?        ��]tc�?��(�"g�?F]t�E�?/�袋.�?�������?�?F]t�E�?]t�E]�?�q�q�?r�q��?      �?      �?              �?      �?      �?      �?                      �?      �?      �?      �?      �?333333�?�������?      �?      �?              �?      �?              �?                      �?      �?                      �?�Mozӛ�?�,d!Y�?a���{�?��=���?;�;��?�؉�؉�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�?�������?      �?        �������?333333�?              �?۶m۶m�?�$I�$I�?�������?�������?UUUUUU�?�������?      �?                      �?      �?      �?              �?      �?              �?        "5�x+��?��sHM0�?9/���?և���X�?              �?      �?      �?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�8��8��?9��8���?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?              �?              �?      �?        9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?�q�q�?�q�q�?              �?      �?        F]t�E�?�.�袋�?              �?UUUUUU�?�������?      �?                      �?���/|*�?�E@V�?              �?GQ栓�?��g|��?+�R��?�	�[���?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �������?�������?;��:���?_�_��?�������?�������?UUUUUU�?UUUUUU�?�������?�������?�q�q�?�q�q�?�������?�������?      �?      �?      �?                      �?      �?              �?                      �?              �?      �?        �z�G��?{�G�z�?���{��?�B!��?              �?�������?�������?      �?        �������?ffffff�?      �?        �?�������?              �?;�;��?ى�؉��?UUUUUU�?UUUUUU�?      �?      �?�������?�������?              �?      �?                      �?      �?        ffffff�?333333�?�$I�$I�?۶m۶m�?F]t�E�?t�E]t�?      �?      �?      �?              �?      �?              �?      �?      �?              �?      �?              �?                      �?      �?        }��|���?���й?�|���?���>��?б�n�Q�?q2�<p�?              �?�1����?�rv��?��N��N�?�؉�؉�?      �?              �?      �?۶m۶m�?�$I�$I�?�$I�$I�?۶m۶m�?      �?      �?333333�?�������?      �?              �?      �?              �?      �?                      �?      �?              �?              �?        �JC��?E'�危?333333�?�����̬?��sHM0�?"5�x+��?�������?UUUUUU�?GX�i���?�{a���?��8��8�?�q�q�?և���X�?9/���?      �?        }g���Q�?W�+�ɕ?      �?              �?      �?      �?      �?              �?      �?              �?        333333�?�������?              �?      �?              �?        �q�q�?�q�q�?      �?      �?      �?                      �?      �?        ]�u]�u�?EQEQ�?      �?        �q�q�?�q�q�?      �?        w�qG�?qG�wĽ?9��8���?�q�q�?۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?      �?      �?���Q��?{�G�z�?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?              �?        �������?�������?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?                      �?      �?      �?      �?                      �??�%C���?�u�y���?              �??���#�?��Gp�?�������?�������?]t�E�?t�E]t�?      �?                      �?L�Ϻ��?к����?      �?      �?t�E]t�?]t�E�?      �?              �?      �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�؉�؉�?;�;��?      �?        �q�q�?�q�q�?      �?                      �?;�;��?;�;��?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?      �?              �?        ��~���?X`��?      �?        �?�?�������?�������?UUUUUU�?UUUUUU�?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ\bshG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                    �?���%&�?�           8�@              O                    �?r�����?U           �@               B                 ��<J@~h����?j             e@              /                    �?     x�?P             `@              .                    �?��
P�?-            �Q@                                  �?:-�.A�?,            �P@                                    @X�Cc�?
             ,@                                   �?r�q��?             @       	       
                 ��@5@      �?             @        ������������������������       �                      @                                hލC@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                  �,@      �?              @        ������������������������       �                      @                                ���,@�q�q�?             @                                 �-@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @               +                    �?r�����?"            �J@                               ���@��k=.��?            �G@        ������������������������       �        	             *@                                 �|Y=@�������?             A@                                  �8@�eP*L��?             &@                                 �5@      �?              @                                   /@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        !       "                 ���4@�㙢�c�?             7@        ������������������������       �                     $@        #       $                 ��2>@�	j*D�?             *@        ������������������������       �                     @        %       *                 `f�A@ףp=
�?             $@        &       '                 X�lA@z�G�z�?             @        ������������������������       �                     @        (       )                    H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ,       -                 �&�)@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        0       5                    �?��o	��?#             M@        1       2                     @ףp=
�?             >@        ������������������������       �                     @        3       4                 ���@�����H�?             ;@        ������������������������       �                     @        ������������������������       �                     8@        6       ?                   `3@؇���X�?             <@       7       8                  ��@�nkK�?             7@        ������������������������       �                      @        9       :                     @��S�ۿ?             .@        ������������������������       �                     �?        ;       >                    �?@4և���?             ,@       <       =                 �|Y=@�C��2(�?	             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        @       A                 03�7@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        C       N                    �?��(\���?             D@       D       G                   �2@$�q-�?            �C@        E       F                 ��e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        H       I                    �?������?             B@       ������������������������       �                     :@        J       K                 p"�X@ףp=
�?             $@       ������������������������       �                     @        L       M                   @E@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        P       �                 03�9@����`�?�            �w@       Q       t                    �?܉���?�            �p@        R       g                    ;@Np�����?#            �I@        S       T                     @l��
I��?             ;@        ������������������������       �                     �?        U       d                    �?�	j*D�?             :@       V       a                   �6@b�2�tk�?
             2@       W       \                   �4@      �?             (@        X       [                    3@�q�q�?             @       Y       Z                 ��!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ]       ^                   �5@X�<ݚ�?             "@        ������������������������       �                      @        _       `                 جJ"@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        b       c                 P�@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        e       f                 P�@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        h       s                    �?      �?             8@       i       j                 ��� @����X�?             5@        ������������������������       �                     @        k       n                 ���&@r�q��?             2@        l       m                   �J@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        o       p                   �A@�8��8��?	             (@       ������������������������       �                     @        q       r                   �C@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        u       �                   �<@��Ujѡ�?�            @k@        v       w                 @3�@����D��?<            @W@       ������������������������       �                     �H@        x       �                   �3@���7�?             F@        y       |                 ��Y @�KM�]�?             3@        z       {                    1@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        }       ~                 ���$@��S�ۿ?
             .@        ������������������������       �                     @               �                   �2@�����H�?             "@        ������������������������       �                     @        �       �                     @r�q��?             @       �       �                   �'@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     9@        �       �                    �?HP�s��?M            @_@       �       �                     �?��ϭ�*�?H             ]@        ������������������������       �                     @        �       �                   @E@�H�@=��?E            �[@       �       �                   @C@���H��?7             U@       �       �                 ��) @����1�?/            @R@       �       �                     @�&=�w��?!            �J@        ������������������������       �                     @        �       �                 �|�>@@9G��?            �H@       �       �                 ��L@ ���J��?            �C@        �       �                 pf�@�����H�?             "@       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     >@        �       �                 �?�@ףp=
�?             $@       ������������������������       �                     @        �       �                   �@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �>@      �?             4@       �       �                     @�n_Y�K�?	             *@        �       �                   �'@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    (@X�<ݚ�?             "@       �       �                 �|�=@�q�q�?             @       �       �                 `��!@���Q��?             @        ������������������������       �                      @        �       �                 ���"@�q�q�?             @        ������������������������       �                     �?        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �D@���!pc�?             &@       �       �                   �C@�<ݚ�?             "@       �       �                     @�q�q�?             @        ������������������������       �                     �?        �       �                 ��	0@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ;@        ������������������������       �                     "@        �       �                    �?2t3����??            �[@        ������������������������       �                    �D@        �       �                 ��$:@��+7��?'            @Q@        ������������������������       �        	             2@        �       �                    D@ҳ�wY;�?            �I@       �       �                   �;@      �?             >@        �       �                    �?      �?              @       �       �                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �>@8�A�0��?             6@        ������������������������       �                     @        �       �                      @     ��?
             0@       �       �                 `f�K@z�G�z�?	             .@       ������������������������       �                     $@        �       �                 �w|c@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?؇���X�?             5@       �       �                    �?ףp=
�?
             4@       �       �                    J@8�Z$���?             *@       �       �                   �G@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                     @�W����?g            �d@       �       �                    N@�Q��k�?5             T@       �       �                   �(@d1<+�C�?2            @R@        ������������������������       �                     �?        �       �                    �?      �?1             R@       �       �                    @�&=�w��?#            �J@        �       �                 ��1V@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        !            �H@        �       �                     �?p�ݯ��?             3@       �       �                   @B@��
ц��?             *@        ������������������������       �                     @        ������������������������       �                     @        �       �                   �3@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �                          @\`*�s�?2             U@       �       �                    �?      �?              H@       �       �                    �?�û��|�?             7@        �       �                   �&@�eP*L��?             &@        ������������������������       �                      @        �       �                 `fV6@�q�q�?             "@       �       �                   �/@؇���X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    )@�q�q�?
             (@        ������������������������       �                     @        �       �                 �y�/@z�G�z�?             @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                       `f7@�J�4�?             9@        �       �                 ��-@�z�G��?             $@        ������������������������       �                     @        �                          �?      �?             @                                 �?���Q��?             @                             �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                              ��T?@��S�ۿ?	             .@       ������������������������       �                     @                                 @      �?              @       	      
                   @r�q��?             @        ������������������������       �                     �?                                �C@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                 @4?,R��?             B@                                �?�>4և��?             <@       ������������������������       �                     &@                                 ,@�t����?             1@                                @z�G�z�?             .@                                @�z�G��?             $@                                @      �?              @        ������������������������       �                     @                                 @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������g *��?�0���M�?��6y_<�?}|�A��?�m۶m��?%I�$I��?     ��?      �?uPuP�?�_�_�?���@���?��~5&�?�m۶m��?%I�$I��?UUUUUU�?�������?      �?      �?              �?      �?      �?      �?                      �?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        Dj��V��?�V�9�&�?g���Q��?br1���?      �?        �������?�������?t�E]t�?]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�7��Mo�?d!Y�B�?      �?        vb'vb'�?;�;��?              �?�������?�������?�������?�������?      �?              �?      �?              �?      �?              �?        �������?UUUUUU�?              �?      �?              �?        ������?���{�?�������?�������?              �?�q�q�?�q�q�?      �?                      �?۶m۶m�?�$I�$I�?�Mozӛ�?d!Y�B�?      �?        �������?�?      �?        n۶m۶�?�$I�$I�?]t�E�?F]t�E�?              �?      �?              �?        �������?333333�?              �?      �?        333333�?�������?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?to��]��?!�8Da�?��k�z�?�Q���?______�?PPPPPP�?Lh/����?h/�����?      �?        vb'vb'�?;�;��?�8��8��?9��8���?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �q�q�?r�q��?              �?�$I�$I�?۶m۶m�?              �?      �?        �������?UUUUUU�?              �?      �?              �?      �?              �?      �?              �?      �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?      �?                      �?              �?��p=�?��A��.�?P?���O�?X`��?      �?        �.�袋�?F]t�E�?�k(���?(�����?      �?      �?      �?                      �?�������?�?      �?        �q�q�?�q�q�?      �?        �������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?              �?        q=
ףp�?{�G�z�?����=�?|a���?      �?        ��+c��?q��$�?�0�0�?��y��y�?�Ν;w��?Ĉ#F��?tHM0���?�x+�R�?      �?        ������?9/���?��-��-�?�A�A�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?;�;��?ى�؉��?      �?      �?      �?                      �?r�q��?�q�q�?UUUUUU�?UUUUUU�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?              �?        F]t�E�?t�E]t�?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?              �?              �?      �?              �?      �?              �?              �?        �}��7��?*A��)�?              �?zӛ����?Y�B��?      �?        �������?�������?      �?      �?      �?      �?      �?      �?      �?                      �?      �?      �?      �?                      �?颋.���?/�袋.�?              �?      �?      �?�������?�������?      �?        �������?333333�?              �?      �?              �?        ۶m۶m�?�$I�$I�?�������?�������?;�;��?;�;��?333333�?�������?      �?                      �?      �?              �?                      �?p>�cp�?��|���?333333�?333333�?�1bĈ�?ݹs�Ν�?      �?              �?      �?�x+�R�?tHM0���?      �?      �?              �?      �?                      �?Cy�5��?^Cy�5�?�؉�؉�?�;�;�?              �?      �?        UUUUUU�?�������?              �?      �?              �?        ��<��<�?b�a��?      �?      �?��,d!�?8��Moz�?]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?      �?                      �?      �?        �z�G��?{�G�z�?ffffff�?333333�?      �?              �?      �?�������?333333�?      �?      �?              �?      �?                      �?      �?        �������?�?      �?              �?      �?�������?UUUUUU�?      �?        �������?�������?              �?      �?              �?        �8��8��?r�q��?�$I�$I�?�m۶m��?      �?        �������?�������?�������?�������?ffffff�?333333�?      �?      �?      �?              �?      �?              �?      �?                      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM!hjh))��}�(h,h/h0M!��h2h3h4hph<�h=Kub������       h                    �?ʡ�;S��?�           8�@               _                    @��6}��?�            �n@              ^                    @$~���?�            �k@              K                 03�5@0@�t�?�            �j@               2                   P,@^����?C            @Z@              %                 `f�%@��+7��?/            @Q@              $                    �?X�Cc�?             E@              #                    �?�	j*D�?            �C@       	       "                 pF%@4�2%ޑ�?            �A@       
                          �1@H�V�e��?             A@        ������������������������       �                     @                                    @      �?             <@        ������������������������       �                      @               !                 X��@@R�}e�.�?             :@                               ��@�+e�X�?             9@                                  �?؇���X�?             ,@                                  �?�C��2(�?             &@        ������������������������       �                      @                                 ��@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                                �|Y:@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                    �?���|���?             &@                               P�N@���Q��?             $@        ������������������������       �                     @                                  �5@؇���X�?             @        ������������������������       �                     @                                pf� @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        &       1                     @�����H�?             ;@       '       (                 `f�)@��2(&�?             6@        ������������������������       �                     @        )       0                    �?     ��?             0@       *       +                    ;@z�G�z�?             .@        ������������������������       �                     �?        ,       -                   �B@؇���X�?             ,@       ������������������������       �                     "@        .       /                    D@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        3       >                    �?X�<ݚ�?             B@        4       9                 ���,@      �?             (@        5       8                    �?���Q��?             @       6       7                   �-@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        :       ;                    �?؇���X�?             @        ������������������������       �                     @        <       =                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ?       H                   @4@�q�q�?             8@       @       A                     @z�G�z�?             4@        ������������������������       �                      @        B       G                    �?�q�q�?             (@       C       D                 �|�;@      �?              @        ������������������������       �                     @        E       F                    .@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        I       J                    ?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        L       ]                    @��Ujѡ�?C            @[@       M       X                    �?X'"7��?B             [@       N       W                 03�<@` A�c̭?;             Y@        O       R                    �?�C��2(�?            �@@        P       Q                    �?      �?             0@        ������������������������       �                      @        ������������������������       �                     ,@        S       T                     @�IєX�?             1@       ������������������������       �        
             .@        U       V                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        (            �P@        Y       Z                     @      �?              @       ������������������������       �                     @        [       \                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        `       a                   -@����X�?             5@        ������������������������       �                     @        b       g                 �|Y:@r�q��?
             2@       c       f                    0@���!pc�?             &@       d       e                 ��T?@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        i                       0�"K@dN�6i��?$           0}@       j                         �B@�ʦ+��?	           �z@       k       �                 `�X.@�ۊ^���?�            �x@       l       {                     @��L��?�            �q@        m       z                    �?���7�?"             F@       n       s                    5@���N8�?!             E@        o       p                   �2@z�G�z�?             @        ������������������������       �                      @        q       r                   �'@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        t       u                   �@@�?�|�?            �B@       ������������������������       �                     9@        v       w                 `f�)@�8��8��?
             (@        ������������������������       �                     @        x       y                   @D@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        |       �                    �?p#�����?�            �m@        }       �                   �6@2L�����?)            @Q@        ~                           �?؇���X�?             @        ������������������������       �                     @        �       �                    -@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��� ��?%             O@       �       �                 �|Y=@Ԫ2��?"            �L@        �       �                  ��@�q�q�?             (@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��S�ۿ?            �F@       �       �                 �|�=@�8��8��?             8@       �       �                 ���@؇���X�?	             ,@        ������������������������       �                     @        �       �                   @@�<ݚ�?             "@       ������������������������       �����X�?             @        ������������������������       �                      @        ������������������������       �                     $@        �       �                 X��A@���N8�?             5@       �       �                  s�@P���Q�?             4@        ������������������������       �                      @        �       �                 ��(@�8��8��?	             (@       ������������������������       �ףp=
�?             $@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?l������?g             e@       �       �                 �?�@�������?d            `d@        �       �                   �7@�}�+r��?1             S@        ������������������������       �                     :@        �       �                   �8@HP�s��?              I@        �       �                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y=@      �?             H@        ������������������������       �        	             *@        �       �                   �@�#-���?            �A@       �       �                 ��@     ��?             0@       ������������������������       �                     (@        �       �                 �&B@      �?             @       �       �                 �|Y>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             3@        �       �                    �?\-��p�?3            �U@       �       �                    �?���O1��?0            �T@       �       �                 @3�@��1��?/            �T@        �       �                    :@�z�G��?             $@        ������������������������       �                     @        �       �                   �A@և���X�?             @       �       �                   �?@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 ���"@�����H�?(             R@       �       �                 0SE @x�}b~|�?             �L@       �       �                   �3@6YE�t�?            �@@        �       �                   �1@      �?             @        ������������������������       �      �?             @        ������������������������       �      �?              @        �       �                 �|�;@�>����?             ;@        ������������������������       �                     $@        �       �                 �|�?@�t����?             1@       �       �                 ��) @z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             8@        �       �                 �|�=@z�G�z�?             .@       �       �                   �<@�8��8��?             (@        ������������������������       �                     @        �       �                 �|Y=@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�c�Α�?E             ]@       �       �                    �?V�a�� �?4            �U@       �       �                    �?����S��?%             M@        �       �                      @�����H�?             "@       �       �                   @@@r�q��?             @        ������������������������       �                     @        �       �                   @G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 `fF:@�J��%�?            �H@        ������������������������       �                     .@        �       �                   �J@��.k���?             A@       �       �                   �<@      �?             8@        ������������������������       �                     @        �       �                 �|�?@�\��N��?
             3@        �       �                   �>@���!pc�?             &@       �       �                 �|Y=@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @G@      �?              @       �       �                   �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 `fF<@ףp=
�?             $@        ������������������������       �                     @        �       �                  )?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?XB���?             =@       ������������������������       �                     9@        �       �                  �v6@      �?             @        ������������������������       �                      @        �       �                 �|�:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?l��[B��?             =@        �       �                 X��@@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          @�û��|�?             7@        �       �                     @���!pc�?             &@        ������������������������       �                     @        �       �                 ��|2@և���X�?             @        ������������������������       �                     @                                  @      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                 �?�8��8��?             (@        ������������������������       �                     @                              �̌4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �@@        	                      03�M@�Gi����?            �B@        
                      03[L@؇���X�?             @                             �|�;@      �?             @        ������������������������       �                      @                              �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �?�z�G��?             >@                                �?      �?             8@                              �̾w@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?                              Ј�U@�n_Y�K�?	             *@       ������������������������       �                     @                              p"�X@      �?              @        ������������������������       �                     @        ������������������������       �                     @                                  �?      �?             @                                �?���Q��?             @                             �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0M!KK��h2h3h4hVh<�h=Kub������������N���I5�?d�~`l��?;ڼOq��?�!XG��?�D�$ �?�������?�Ե���?Ċ����?�K��K��?6Z�5Z��?Y�B��?zӛ����?�m۶m��?%I�$I��?;�;��?vb'vb'�?�A�A�?�������?ZZZZZZ�?iiiiii�?              �?      �?      �?              �?�;�;�?'vb'vb�?���Q��?R���Q�?�$I�$I�?۶m۶m�?F]t�E�?]t�E�?              �?�q�q�?�q�q�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?]t�E]�?�������?333333�?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?      �?              �?              �?              �?        �q�q�?�q�q�?t�E]t�?��.���?              �?      �?      �?�������?�������?      �?        �$I�$I�?۶m۶m�?              �?�������?333333�?      �?                      �?              �?              �?�q�q�?r�q��?      �?      �?333333�?�������?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        �������?�������?      �?                      �?              �?      �?      �?      �?                      �?��A��.�?��p=�?B{	�%��?Lh/����?���Q��?
ףp=
�?F]t�E�?]t�E�?      �?      �?      �?                      �?�?�?              �?      �?      �?              �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?                      �?              �?      �?        ���u�a�?0��(�y�?'9�t��?c?-���?���x��?Z�����?����?�\���?�.�袋�?F]t�E�?��y��y�?�a�a�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        *�Y7�"�?к����?      �?        UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?        7a~W��?�#{���?�k�ځ�?�Q�g���?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        �{����?�B!��?$���>��?p�}��?�������?�������?      �?                      �?�������?�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        9��8���?�q�q�?�m۶m��?�$I�$I�?      �?              �?        ��y��y�?�a�a�?ffffff�?�������?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?              �?              �?        �a�a�?=��<��?��Ŗ���?)��I� �?�5��P�?(�����?      �?        q=
ףp�?{�G�z�?      �?      �?      �?                      �?      �?      �?      �?        �A�A�?_�_�?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        a����?�{a���?P�M�_�?���ˊ��?�+Q���?,Q��+�?ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?        �q�q�?�q�q�?�YLg1�?Lg1��t�?'�l��&�?e�M6�d�?      �?      �?      �?      �?      �?      �?�Kh/��?h/�����?      �?        <<<<<<�?�?�������?�������?      �?                      �?      �?              �?        �������?�������?UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?333333�?              �?      �?        5�rO#,�?�{a���?��{a�?a���{�?X�i���?O#,�4��?�q�q�?�q�q�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        c}h���?9/����?      �?        �������?�?      �?      �?              �?�5��P�?y�5���?F]t�E�?t�E]t�?�������?333333�?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        GX�i���?�{a���?      �?              �?      �?      �?              �?      �?      �?                      �?���=��?GX�i���?UUUUUU�?�������?              �?      �?        8��Moz�?��,d!�?t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?              �?      �?              �?        o0E>��?#�u�)��?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?                      �?              �?ffffff�?333333�?      �?      �?]t�E�?F]t�E�?      �?                      �?;�;��?ى�؉��?      �?              �?      �?              �?      �?              �?      �?333333�?�������?      �?      �?              �?      �?                      �?              �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJj�c;hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       P                    �?|��;;��?�           8�@               O                    @� ��1�?�            �n@                                  �?�+$�jP�?�            `n@                                   @�<p���?4            �T@                                   @p=
ףp�?3             T@       ������������������������       �                    �E@                                  �,@��G���?            �B@        ������������������������       �                     @        	                           �?��a�n`�?             ?@        
                        `�@1@      �?	             (@                                  �?�q�q�?             "@                                 �7@      �?             @        ������������������������       �                     �?                                   �?�q�q�?             @        ������������������������       �                     �?                                �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �-@z�G�z�?             @        ������������������������       �                      @                                �|Y6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                ���@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                      @               0                     @�_�8�?j             d@              -                 ���a@ ���v��?B            �X@              *                   �K@�zvܰ?;             V@               )                   �+@ Df@��?8            �T@        !       "                   �'@�C��2(�?             6@        ������������������������       �                     &@        #       (                   �B@"pc�
�?             &@       $       '                    ;@ףp=
�?             $@        %       &                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        )            �N@        +       ,                 `f�2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        .       /                 03c@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        1       F                 ���1@      �?(             O@       2       =                 P��%@��]�T��?            �D@       3       <                   �"@8�A�0��?             6@       4       ;                    �?     ��?             0@       5       :                    �?��
ц��?
             *@       6       9                    ;@�q�q�?	             (@       7       8                 xF� @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        >       E                    �?�KM�]�?             3@       ?       @                    �?�t����?
             1@        ������������������������       �                      @        A       B                 P��)@�<ݚ�?             "@        ������������������������       �                      @        C       D                 �|�<@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        G       N                    @���N8�?             5@       H       M                 �̼6@�S����?             3@        I       J                 03C3@      �?              @        ������������������������       �                     @        K       L                     @���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     @        Q       d                    @� j����?            }@        R       S                 @3�4@�t����?             1@        ������������������������       �                     @        T       _                    @�eP*L��?
             &@       U       V                    �?և���X�?             @        ������������������������       �                     �?        W       \                    �?�q�q�?             @       X       [                   l@@      �?             @       Y       Z                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ]       ^                 pf�X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        `       c                 ��T?@      �?             @        a       b                 03�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        e       �                     �?���X�?            |@        f       �                 �̾w@�^�X�?<            @X@       g       r                   �<@��n%�4�?:            �W@        h       o                    �?      �?             0@       i       j                 ���Q@�z�G��?	             $@       ������������������������       �                     @        k       n                  "&d@      �?             @        l       m                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        p       q                    7@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        s       �                   @@@����?.            �S@        t       �                    �?ȵHPS!�?             :@       u       z                    �?�LQ�1	�?             7@        v       w                 ���<@�����H�?             "@        ������������������������       �                     @        x       y                 03SA@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        {       �                   �>@؇���X�?             ,@        |       }                 `fF<@����X�?             @       ������������������������       �                     @        ~                        �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�	j*D�?             J@       �       �                    @@z�G�z�?            �A@       �       �                 ���=@�q�q�?             5@       �       �                    �?�<ݚ�?             2@       �       �                    �?      �?
             0@        ������������������������       �                      @        �       �                 ��I*@����X�?	             ,@        ������������������������       �                     @        �       �                    D@���|���?             &@        ������������������������       �                      @        �       �                 `f�;@�<ݚ�?             "@       �       �                   �J@����X�?             @        �       �                    H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     ,@        �       �                 `�iJ@��.k���?             1@        ������������������������       �                     @        �       �                 `ށK@և���X�?             ,@        ������������������������       �                      @        �       �                 ЈT@      �?             (@        ������������������������       �                     @        �       �                    �?�q�q�?             "@        ������������������������       �                     @        �       �                   �D@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �                          @Ha�>i�?�            �u@       �                       �̄H@L��rH�?�            Pu@       �       �                    ,@l������?�             u@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �                          �?������?�            �t@       �                         �*@0D#��^�?�            �q@       �       �                    �?�K��G^�?�            @p@        �       �                     @r�q��?!             K@        ������������������������       �                      @        �       �                    �?D>�Q�?             J@       �       �                 ���@r�q��?             >@        �       �                 03S@@4և���?             ,@        ������������������������       �                     @        �       �                 �|�9@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y=@      �?	             0@        ������������������������       �                     @        ������������������������       �                     (@        �       �                 �|Y=@"pc�
�?             6@        ������������������������       �                      @        �       �                 ���@ףp=
�?             4@        ������������������������       �                     @        �       �                 X��A@؇���X�?	             ,@       �       �                 ��(@r�q��?             (@       ������������������������       �z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                 �?�@\�t��Y�?|            �i@        �       �                 �Yu@,N�_� �?1            �R@       �       �                    7@`�H�/��?             �I@        ������������������������       �                     7@        �       �                 ��L@�>4և��?             <@       �       �                 �|Y>@ȵHPS!�?             :@       �       �                 �&b@@�0�!��?             1@        ������������������������       �                     @        �       �                 ���@      �?             (@        ������������������������       �                     �?        �       �                 �|Y;@"pc�
�?             &@       ������������������������       �                     @        �       �                 ��,@����X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     7@        �       �                   �:@�禺f��?K            �`@        �       �                     @`Ӹ����?            �F@        �       �                    5@$�q-�?             *@        �       �                    &@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 pf� @      �?             @@        �       �                 @3�@@4և���?	             ,@        ������������������������       �                     @        �       �                   �1@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        
             2@        �       �                 @3�@�����?-            �U@        �       �                   �?@      �?              @        ������������������������       �                     @        �       �                   �A@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                   �;@��r�Z}�?)            �S@        �       �                 ���%@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��) @�?�'�@�?'             S@        ������������������������       �                     7@        �       �                     @r�����?            �J@       �       �                   �F@�����H�?             B@       �       �                 `fF)@"pc�
�?             6@        ������������������������       �                     @        �       �                    @@������?             1@        ������������������������       �                     "@        �       �                   @B@      �?              @        ������������������������       �                     @        �       �                   @D@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     ,@        �       �                 pF� @ҳ�wY;�?	             1@        ������������������������       �                      @        �       �                 ���"@������?             .@        ������������������������       �                      @        �       �                   �<@և���X�?             @        ������������������������       �                     �?        �                        �|Y=@�q�q�?             @        ������������������������       �                     @                              �|�=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@                                 �? "��u�?!             I@                              03�-@؇���X�?             5@        ������������������������       �                     @              	                ��.@z�G�z�?	             .@        ������������������������       �                     �?        
                         �?؇���X�?             ,@                                �?�8��8��?             (@        ������������������������       �                     @                                 �?r�q��?             @                                 @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                               �v6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     =@                                 >@���Q��?             @                                ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������|d�_Z�?�7s@K�?������?������?B{	�%��?/�����?�����?}���|�?ffffff�?333333�?              �?v�)�Y7�?#�u�)��?              �?�s�9��?�c�1��?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?(�����?�5��P�?      �?                      �?      �?        �O���? l<�?��?1ogH�۩?�y;Cb�?t�E]t�?颋.���?��k���?c��7�:�?F]t�E�?]t�E�?              �?F]t�E�?/�袋.�?�������?�������?      �?      �?      �?                      �?              �?      �?                      �?�������?�������?      �?                      �?F]t�E�?/�袋.�?      �?                      �?      �?      �?jW�v%j�?KԮD�J�?颋.���?/�袋.�?      �?      �?�;�;�?�؉�؉�?�������?�������?UUUUUU�?�������?              �?      �?              �?                      �?              �?      �?        (�����?�k(���?�?<<<<<<�?              �?�q�q�?9��8���?              �?�$I�$I�?�m۶m��?      �?                      �?              �?�a�a�?��y��y�?(������?^Cy�5�?      �?      �?      �?        �������?333333�?              �?      �?              �?                      �?      �?        JZ���I�?ٖ�m���?�������?�������?              �?]t�E�?t�E]t�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?              �?              �?      �?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?۶m۶��?�$I�$I�?���Id�?��4l7��?������?���
b�?      �?      �?333333�?ffffff�?              �?      �?      �?      �?      �?      �?                      �?      �?        �������?UUUUUU�?      �?                      �?H�4H�4�?��-��-�?��N��N�?�؉�؉�?��Moz��?Y�B��?�q�q�?�q�q�?      �?        �������?�������?              �?      �?        ۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        vb'vb'�?;�;��?�������?�������?UUUUUU�?UUUUUU�?9��8���?�q�q�?      �?      �?      �?        �m۶m��?�$I�$I�?      �?        ]t�E]�?F]t�E�?              �?9��8���?�q�q�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?                      �?      �?        �?�������?              �?�$I�$I�?۶m۶m�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?2��C�?sޑ�3�?'�p�	'�?�{�Ǿ?�a�a�?=��<��?UUUUUU�?UUUUUU�?      �?                      �?��g�`��?к����?G#ƿD�?��&�ڽ??�?��?�?�?�?�������?UUUUUU�?      �?        b'vb'v�?vb'vb'�?�������?UUUUUU�?n۶m۶�?�$I�$I�?      �?              �?      �?              �?      �?              �?      �?              �?      �?        /�袋.�?F]t�E�?              �?�������?�������?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?�������?�������?      �?              �?        P ���E�?��VCӽ?h�`�|��?���L�?�������?�?      �?        �$I�$I�?�m۶m��?��N��N�?�؉�؉�?ZZZZZZ�?�������?      �?              �?      �?              �?/�袋.�?F]t�E�?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        e�M6�d�?m��&�l�??�>��?l�l��?�؉�؉�?;�;��?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?              �?      �?n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?        ;���C��?/�I��?      �?      �?              �?333333�?�������?      �?      �?      �?        G�D�#�?�&��jq�?UUUUUU�?UUUUUU�?              �?      �?        ������?y�5���?      �?        Dj��V��?�V�9�&�?�q�q�?�q�q�?/�袋.�?F]t�E�?      �?        xxxxxx�?�?      �?              �?      �?              �?�������?�������?      �?              �?      �?      �?        �������?�������?              �?wwwwww�?�?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �G�z�?���Q��?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJGԙGhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMMhjh))��}�(h,h/h0MM��h2h3h4hph<�h=Kub������       �                     @e�L��?�           8�@               o                   �D@.������?�            �t@                                  �?t�C�#��?�            �m@                                   �?���#�İ?C            �]@                                  �?�k~X��?'             R@        ������������������������       �                     3@                                  �+@�O4R���?            �J@                                  �9@`2U0*��?             9@        	       
                   �'@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     <@                                ���a@���.�6�?             G@                                   �? qP��B�?            �E@        ������������������������       �                     3@                                   �? �q�q�?             8@        ������������������������       �                     @                                   6@�}�+r��?             3@                                  �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             1@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               N                     �?�0�w�?Q            �]@               5                    �?:2vz�M�?(            �N@               4                 �̾w@��S���?             >@              3                 �U�X@�5��?             ;@              .                   �A@      �?             6@               #                   �8@�q�q�?             .@        !       "                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        $       -                    �?      �?	             (@       %       &                 �|Y<@      �?              @        ������������������������       �                      @        '       ,                   @@@      �?             @       (       +                 ��2>@      �?             @        )       *                 ���<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        /       2                    �?؇���X�?             @       0       1                    C@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        6       7                 03:@���@M^�?             ?@        ������������������������       �                     "@        8       I                    �?�eP*L��?             6@       9       H                    �?��.k���?             1@       :       E                   �>@     ��?             0@        ;       <                 03k:@z�G�z�?             $@        ������������������������       �                     @        =       D                   @>@����X�?             @       >       ?                 �|Y=@�q�q�?             @        ������������������������       �                     �?        @       C                 `fF<@z�G�z�?             @       A       B                 �|�?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        F       G                 �|�<@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        J       K                    <@���Q��?             @        ������������������������       �                      @        L       M                 03�S@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        O       f                    �?д>��C�?)             M@       P       e                 ���?@���H��?             E@       Q       X                   �)@��(\���?             D@       R       S                    �?�nkK�?             7@        ������������������������       �                      @        T       W                    5@���N8�?             5@        U       V                    &@؇���X�?             @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     ,@        Y       Z                    �?�t����?             1@        ������������������������       �                     �?        [       \                 �|Y<@      �?             0@        ������������������������       �                      @        ]       ^                 �|�=@      �?              @        ������������������������       �                     �?        _       d                   �3@؇���X�?             @       `       a                    @@r�q��?             @        ������������������������       �                      @        b       c                   �A@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        g       h                    �?     ��?             0@        ������������������������       �                      @        i       j                   @.@      �?              @        ������������������������       �                     �?        k       l                    :@����X�?             @        ������������������������       �                     @        m       n                    0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        p       }                    �?VP��g��?:             W@        q       z                     �?"pc�
�?             6@       r       y                   �I@�C��2(�?
             &@        s       x                    �?      �?             @       t       u                 0#R;@�q�q�?             @        ������������������������       �                     �?        v       w                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        {       |                   �K@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ~       �                   �J@������?+            �Q@              �                 `ff:@RB)��.�?            �E@        ������������������������       �        	             3@        �       �                 `f�:@      �?             8@        �       �                   @G@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        �       �                    �?�<ݚ�?             2@       �       �                 0��M@@�0�!��?             1@       �       �                    �?���!pc�?	             &@        ������������������������       �                     �?        �       �                    �?z�G�z�?             $@        �       �                   @A@z�G�z�?             @        �       �                   �=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     �?z�G�z�?             @       �       �                    G@      �?             @       �       �                  x#J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ;@        �       �                    �?:��r:�?�            �w@        �       �                    �?������?E            �[@        �       �                 X�,A@      �?             @@       �       �                 P��+@д>��C�?             =@       �       �                    �?�IєX�?             1@        ������������������������       �                     @        �       �                 �|�9@$�q-�?	             *@        ������������������������       �                      @        �       �                 ���@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?�q�q�?
             (@       �       �                    �?      �?              @       �       �                    @և���X�?             @       �       �                 �|�7@�q�q�?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                 P�h2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��i @p`q�q��?-            �S@       �       �                 �|Y=@�U�:��?!            �M@        �       �                    �?      �?              @       �       �                    �?����X�?             @       �       �                   @9@      �?             @        ������������������������       �                      @        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                  ��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �I@        �       �                    �?�G�z��?             4@       �       �                 ��$1@���|���?             &@        ������������������������       �                     @        �       �                   �2@      �?              @        ������������������������       �                     @        �       �                 03�7@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       L                   @��0p'��?�            �p@       �                          �?�����?�            Pp@       �                       ��C@��v����?�             i@       �       �                    �?<$c*(��?}            `h@        �       �                   �6@���!pc�?            �@@        �       �                    �?�eP*L��?	             &@       �       �                 ���@�q�q�?             "@        ������������������������       �                     @        �       �                    '@      �?             @        ������������������������       �                     �?        �       �                  �#@���Q��?             @       �       �                    4@      �?             @        ������������������������       �                      @        �       �                 �̜!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �&B@��2(&�?             6@        ������������������������       �                     @        �       �                     @r�q��?
             2@       �       �                   �9@�t����?	             1@        ������������������������       �                     @        �       �                    �?"pc�
�?             &@       �       �                  SE"@      �?              @       �       �                 P��@�q�q�?             @        ������������������������       �                     �?        �       �                 ��� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �                         �<@ wVX(6�?h            @d@       �       �                    �?(�5�f��?5            �S@       �       �                   �0@��.N"Ҭ?.            @Q@        �       �                 pFD!@؇���X�?             @       �       �                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        �       �                   �:@0�z��?�?)             O@       ������������������������       �        !             I@        �       �                 �� @�8��8��?             (@       ������������������������       �                      @        �       �                   �;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 P�@ףp=
�?             $@       ������������������������       �                     @        �       �                    2@�q�q�?             @        ������������������������       �                     �?        �                           �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?�o��gn�?3            �T@                               @@@�ӭ�a��?,             R@                             �|�=@��[�8��?            �I@             
                ��) @�ݜ�?            �C@             	                 sW@�g�y��?             ?@                              pf�@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@                              pf� @      �?              @        ������������������������       �                      @                              ���"@�q�q�?             @        ������������������������       �                     @                              �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                �?@      �?             (@                             �?�@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                              P�@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     5@        ������������������������       �                     &@                                 ;@�q�q�?             @        ������������������������       �                     @                              �|�>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?               /                   �?���Q��?)             N@        !      (                   �?����X�?
             ,@       "      '                   @�<ݚ�?             "@       #      &                   ,@      �?              @        $      %                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        )      ,                   �?���Q��?             @        *      +                @3�,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        -      .                  �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        0      =                   @8����?             G@        1      4                   �?���Q��?
             .@        2      3                ��|2@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        5      8                   @      �?              @        6      7                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        9      :                   �?z�G�z�?             @        ������������������������       �                      @        ;      <                ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        >      K                   �?�חF�P�?             ?@       ?      H                   �?�E��ӭ�?             2@       @      E                   @      �?              @       A      B                `fv1@z�G�z�?             @        ������������������������       �                      @        C      D                ���5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        F      G                   @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        I      J                   ,@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     $@        �*       h�h))��}�(h,h/h0MMKK��h2h3h4hVh<�h=Kub������������v�S(��?��X��?�q���?3� ?7�?��7a~�?��td�@�?'u_[�?��N��?�q�q�?�8��8��?              �?�x+�R�?:�&oe�?{�G�z�?���Q��?      �?      �?              �?      �?                      �?              �?Y�B��?���7���?�}A_З?��}A�?              �?UUUUUU�?�������?              �?(�����?�5��P�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        v�Qv�Q�?�\�\�?��6�S\�?��!XG�?�?�������?h/�����?/�����?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?              �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?              �?                      �?�s�9��?�c�1��?      �?        ]t�E�?t�E]t�?�?�������?      �?      �?�������?�������?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�������?UUUUUU�?              �?      �?              �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?a���{�?|a���?�0�0�?��y��y�?�������?333333�?�Mozӛ�?d!Y�B�?      �?        ��y��y�?�a�a�?۶m۶m�?�$I�$I�?      �?      �?      �?              �?        <<<<<<�?�?      �?              �?      �?      �?              �?      �?              �?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?              �?                      �?      �?      �?      �?              �?      �?      �?        �$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?        �Mozӛ�?-d!Y��?F]t�E�?/�袋.�?F]t�E�?]t�E�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?              �?t�E]t�?F]t�E�?              �?      �?        ,��+���?PuPu�?S֔5eM�?���)k��?      �?              �?      �?UUUUUU�?�������?      �?      �?              �?9��8���?�q�q�?ZZZZZZ�?�������?F]t�E�?t�E]t�?              �?�������?�������?�������?�������?      �?      �?      �?                      �?      �?        �������?�������?      �?      �?      �?      �?      �?                      �?      �?              �?              �?                      �?      �?        �i���`�?vX�Q�}�?G���w�?q��$�?      �?      �?|a���?a���{�?�?�?              �?;�;��?�؉�؉�?              �?F]t�E�?]t�E�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?      �?        
�Z܄�?�3����?�A�I�?�pR�屵?      �?      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?]t�E]�?F]t�E�?      �?              �?      �?      �?        �������?�������?              �?      �?        �q�q�?9��8���?              �?      �?        �&�U��?e��?;���C��?/�I��?5&����?*g��1�?��9��9�?�1�1�?F]t�E�?t�E]t�?]t�E�?t�E]t�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?333333�?�������?      �?      �?      �?              �?      �?              �?      �?                      �?      �?        ��.���?t�E]t�?      �?        �������?UUUUUU�?<<<<<<�?�?      �?        /�袋.�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?                      �?k~X�<�?�<ݚ�?�=Q���?�&��jq�?�3J���?ہ�v`��?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        |���{�?�B!��?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        rY1P��?�7�:���?�q�q�?�8��8��?�?�������?\��[���?�i�i�?��{���?�B!��?�q�q�?�q�q�?      �?                      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?۶m۶m�?�$I�$I�?      �?                      �?333333�?�������?              �?      �?      �?      �?              �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?�$I�$I�?�m۶m��?�q�q�?9��8���?      �?      �?      �?      �?              �?      �?                      �?      �?        �������?333333�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        d!Y�B�?8��Moz�?�������?333333�?۶m۶m�?�$I�$I�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�Zk����?��RJ)��?�q�q�?r�q��?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��AhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       V                    �?�4�O��?�           8�@               ;                    �?��%�[H�?�            `o@              0                  S�-@�nW��?{            @i@                                    @��]�T��?6            �T@                                   �?z�G�z�?             9@        ������������������������       �                     @               
                   �'@�d�����?             3@              	                   �J@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @                                   B@      �?              @       ������������������������       �                     @                                   D@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @               )                 �|�<@T�7�s��?&            �L@                                  �?�Gi����?            �B@                                   �?"pc�
�?             &@                                 �,@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @               &                    �?�θ�?             :@              #                    �?��<b���?             7@                                  3@������?             1@                                P��@�q�q�?             @        ������������������������       �                     �?                                ��!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               "                   �7@؇���X�?             ,@               !                 pff@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        $       %                    4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        '       (                    -@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        *       /                 ���*@R���Q�?             4@       +       ,                    �?�KM�]�?             3@       ������������������������       �        	             *@        -       .                 ��� @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        1       :                    @��(\���?E             ^@       2       3                    �?���͡?A            @\@        ������������������������       �                     I@        4       5                     �?�i�y�?$            �O@        ������������������������       �                     ;@        6       9                    �?�X�<ݺ?             B@       7       8                   �E@�>����?             ;@       ������������������������       �                     9@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        <       M                    @ڡR����?"            �H@       =       L                    @��
P��?            �A@       >       C                    �?     ��?             @@        ?       @                     @      �?             $@        ������������������������       �                     @        A       B                 �|Y=@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        D       I                     @8�A�0��?             6@       E       H                     �?z�G�z�?             .@        F       G                    )@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        J       K                 @34@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        N       U                 �|Y7@؇���X�?             ,@       O       P                 ���3@�<ݚ�?             "@        ������������������������       �                     �?        Q       T                    @      �?              @        R       S                    @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        W       �                   �/@>W]���?           �|@       X       Y                 ���@�yL�x��?�            �r@        ������������������������       �                     @@        Z       [                    ,@ �Zz�q�?�            �p@        ������������������������       �                      @        \       �                   @E@�~�H��?�            pp@       ]       �                   �D@ �����?�             m@       ^       _                 ��@h�˹�?�            �l@        ������������������������       �                      @        `       �                   �?@ ڀ��/�?�            @l@       a       ~                 @3�@��a�n`�?t            @g@        b       }                    �?��S�ۿ?7            �V@       c       |                 �?$@���M�?6            @V@       d       e                 ���@�q��/��?            �H@        ������������������������       �                     @        f       u                    �?؇���X�?             E@       g       h                   �5@�GN�z�?             6@        ������������������������       �                      @        i       t                    �?R���Q�?             4@       j       q                  s�@r�q��?             2@       k       p                 `��@�C��2(�?             &@       l       m                 �|=@      �?              @        ������������������������       �                      @        n       o                 �|�=@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     @        r       s                 �|Y=@����X�?             @        ������������������������       �                     �?        ������������������������       �r�q��?             @        ������������������������       �                      @        v       w                 �|�;@P���Q�?             4@       ������������������������       �                     .@        x       y                 ��,@z�G�z�?             @        ������������������������       �                      @        z       {                 �|Y>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     D@        ������������������������       �                     �?               �                    �?      �?=             X@       �       �                     @d۬����?;            @W@        �       �                    4@$�q-�?             :@        �       �                   �2@�q�q�?             @        ������������������������       �                      @        �       �                   �'@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     4@        �       �                    �?��v����?*            �P@       �       �                   �0@R���Q�?'             N@        �       �                 pFD!@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 `�X#@X�;�^o�?$            �K@       �       �                   �:@؇���X�?             �H@       �       �                   �3@�>����?             ;@        �       �                   �1@"pc�
�?             &@        ������������������������       �                     @        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        �       �                 0S5 @z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                    �?�GN�z�?             6@        ������������������������       �                      @        �       �                 ��) @      �?             4@       ������������������������       �                     (@        �       �                 pf� @      �?              @        ������������������������       �                     �?        �       �                   �;@և���X�?             @        ������������������������       �                      @        �       �                 ��)"@���Q��?             @        ������������������������       �                     �?        �       �                   �<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��*@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @A@z�G�z�?             D@        �       �                    �?�����?             3@       �       �                 `fF)@�q�q�?             2@       �       �                    �?8�Z$���?	             *@        ������������������������       �                     @        �       �                   @@@z�G�z�?             $@        �       �                   �@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �@@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @C@���N8�?             5@       ������������������������       �                     (@        �       �                    �?�����H�?             "@       �       �                 �?�@؇���X�?             @        ������������������������       �                     @        �       �                     @�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                     @���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     >@        �       �                     �?��0�=8�?a            `d@        �       �                  �>@T�iA�?,            �Q@        �       �                   �F@�d�����?             3@       ������������������������       �                      @        �       �                   @=@�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�t����?!            �I@       �       �                    �?�'�`d�?            �@@        �       �                   �7@      �?
             0@        ������������������������       �                     @        �       �                 �̾w@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        �       �                 `��S@@�0�!��?
             1@       ������������������������       �                     *@        �       �                 �|�0@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?X�<ݚ�?             2@       �       �                   �G@���|���?
             &@       �       �                    C@      �?              @       �       �                    �?�q�q�?             @        �       �                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    =@      �?             @        ������������������������       �                     �?        �       �                   @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��f`@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �                           �?��a�n`�?5            @W@        �       �                    �?>A�F<�?             C@        �       �                    �?���|���?             &@       �       �                 ��d5@      �?              @        �       �                   �2@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 03�7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    9@�����H�?             ;@        ������������������������       �                      @        �       �                     @�S����?             3@        ������������������������       �                     "@        �       �                    �?�z�G��?             $@        �       �                 �|�;@���Q��?             @        ������������������������       �                      @        �       �                 �|�>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 @^(��I�?            �K@                             03{3@h+�v:�?             A@                                �:@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                 :@����X�?             <@                             03c4@b�2�tk�?             2@        ������������������������       �                     @        	      
                �̌4@��
ц��?             *@        ������������������������       �                     @                              ��\6@���Q��?             $@                                 +@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 �?�q�q�?             @        ������������������������       �                     @                                �3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?                                 �?���N8�?             5@       ������������������������       �                     *@                              pf�C@      �?              @                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������X�>�?2�N����?D�Tw�V�?^�UD�T�?�y��~��?��Q`��?jW�v%j�?KԮD�J�?�������?�������?              �?y�5���?Cy�5��?F]t�E�?/�袋.�?              �?      �?              �?      �?              �?333333�?�������?      �?                      �?�}��?p�}��?o0E>��?#�u�)��?F]t�E�?/�袋.�?�$I�$I�?�m۶m��?              �?      �?                      �?ى�؉��?�؉�؉�?��,d!�?��Moz��?xxxxxx�?�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        �������?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        333333�?333333�?(�����?�k(���?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        333333�?�������?x�!���?$��Co�?              �?AA�?�������?              �?�q�q�?��8��8�?h/�����?�Kh/��?              �?      �?                      �?      �?        ����S��?����X�?_�_��?PuPu�?      �?      �?      �?      �?              �?�������?UUUUUU�?              �?      �?        /�袋.�?颋.���?�������?�������?۶m۶m�?�$I�$I�?      �?                      �?              �?۶m۶m�?�$I�$I�?              �?      �?              �?        ۶m۶m�?�$I�$I�?9��8���?�q�q�?              �?      �?      �?      �?      �?      �?                      �?      �?              �?        &��~]�?i��s��?��X��?*7�9u��?      �?        Γ�ȰA�?�a��y�?              �?�H�x�?���-g:�?)#�e�?���X�ܿ?^Cy�5�?�5��P�?              �?�\�(�u�?�Ź�Q�?�s�9��?�c�1Ƹ?�������?�?��^����?�E(B�?/����?և���X�?      �?        ۶m۶m�?�$I�$I�?�袋.��?]t�E�?              �?333333�?333333�?�������?UUUUUU�?]t�E�?F]t�E�?      �?      �?      �?        �������?UUUUUU�?      �?      �?      �?              �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        ffffff�?�������?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?      �?7�p�7�?Hy�G�?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        5&����?*g��1�?333333�?333333�?333333�?�������?              �?      �?        �־a��?J��yJ�?۶m۶m�?�$I�$I�?�Kh/��?h/�����?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?      �?              �?        �袋.��?]t�E�?      �?              �?      �?      �?              �?      �?              �?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?              �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?ffffff�?ffffff�?Q^Cy��?^Cy�5�?UUUUUU�?UUUUUU�?;�;��?;�;��?      �?        �������?�������?      �?      �?              �?      �?              �?        �������?�������?      �?                      �?      �?        ��y��y�?�a�a�?      �?        �q�q�?�q�q�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        333333�?�������?UUUUUU�?UUUUUU�?      �?              �?        �g*�/�?�0�Qġ�?�+��+��?;��:���?y�5���?Cy�5��?              �?]t�E�?t�E]t�?      �?                      �?�������?�������?6�d�M6�?'�l��&�?      �?      �?              �?�؉�؉�?;�;��?      �?                      �?ZZZZZZ�?�������?      �?              �?      �?              �?      �?        r�q��?�q�q�?F]t�E�?]t�E]�?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?�c�1��?�s�9��?������?Cy�5��?]t�E]�?F]t�E�?      �?      �?333333�?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?      �?        (������?^Cy�5�?      �?        ffffff�?333333�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �7�}���?J��yJ�?�������?xxxxxx�?UUUUUU�?�������?              �?      �?        �m۶m��?�$I�$I�?�8��8��?9��8���?      �?        �؉�؉�?�;�;�?              �?333333�?�������?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?                      �?��y��y�?�a�a�?      �?              �?      �?      �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ,�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������       d                     @>AU`�z�?�           8�@               ;                     �?���H.�?�            �r@              :                    @��$
���?m            `c@                                  �?ҳ�wY;�?l             c@                                   "@ �й���?0            @R@        ������������������������       �                     �?        ������������������������       �        /             R@                                 �>@��Q���?<             T@        	                          @L@      �?             8@       
                        03:@�X����?             6@        ������������������������       �                     @                                   @@r�q��?             2@                                �|�=@�z�G��?             $@                                  �?      �?              @                                �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @               3                    �?d}h���?+             L@              $                    �?�5��
J�?$             G@              #                 p�w@ȵHPS!�?             :@              "                    �?HP�s��?             9@                                �|Y<@"pc�
�?
             &@                                 �}S@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               !                 p�i@@�����H�?             "@                                  �>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     �?        %       (                    =@���Q��?             4@        &       '                 �U�X@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        )       *                 �5L@������?             .@        ������������������������       �                     @        +       0                   �G@���|���?             &@        ,       -                 03�U@r�q��?             @        ������������������������       �                     @        .       /                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       2                 @�pX@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        4       9                    �?ףp=
�?             $@       5       6                    �?�����H�?             "@       ������������������������       �                     @        7       8                  "&d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        <       _                    �?l��[B��?Z             b@       =       ^                   �E@�	j*D�?>            �V@       >       ?                    @:%�[��?3            �Q@        ������������������������       �                     @        @       S                    �?�萻/#�?0            �P@        A       L                    �? �Cc}�?             <@       B       C                    �?�KM�]�?             3@        ������������������������       �                     @        D       K                   �B@؇���X�?             ,@       E       F                 `f�)@$�q-�?             *@        ������������������������       �                     @        G       J                    1@�����H�?             "@       H       I                    ;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        M       N                   �9@�����H�?             "@        ������������������������       �                     @        O       R                   �7@z�G�z�?             @        P       Q                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       ]                 �|�=@$�q-�?            �C@       U       \                   �3@H%u��?             9@       V       [                 �|�<@r�q��?
             2@       W       Z                    &@      �?	             0@        X       Y                   �7@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     4@        `       a                    <@H�ՠ&��?             K@       ������������������������       �                     B@        b       c                    �?b�2�tk�?	             2@       ������������������������       �                     &@        ������������������������       �                     @        e       �                    @,�+Ά1�?�            �y@       f       �                 `�X.@&�
�M�?�            �w@       g       ~                    �?ܱ#_��?�            `r@        h       }                    A@��h!��?#            �L@       i       z                    �? s�n_Y�?             J@       j       q                 �̌@��0{9�?            �G@       k       l                 �|�;@�IєX�?             A@        ������������������������       �                     &@        m       p                 ���@���}<S�?             7@        n       o                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             2@        r       s                    �?�n_Y�K�?	             *@        ������������������������       �                     @        t       y                    �?X�<ݚ�?             "@       u       x                 ��� @�q�q�?             @       v       w                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        {       |                    .@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               �                    �?�BѶ�n�?�            �m@       �       �                 ���@X�M|H�?�            `k@        ������������������������       �                     1@        �       �                 ��@��x��?s            @i@        ������������������������       �                     �?        �       �                   �0@�qM�R��?r             i@        �       �                    �?�q�q�?             @       �       �                 pf�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�"P��?o            �h@        �       �                 �|Y=@x�����?            �C@        �       �                    ;@և���X�?             @       �       �                 ��@      �?             @       �       �                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��(@      �?             @@       �       �                 �|�=@"pc�
�?             6@       �       �                 ���@������?
             1@        ������������������������       �                     @        �       �                    �?����X�?             ,@        ������������������������       �                     �?        �       �                 �Y�@�θ�?             *@        ������������������������       �                     �?        ������������������������       �      �?             (@        ������������������������       �                     @        ������������������������       �                     $@        �       �                 �?�@�<� w�?V            �c@       �       �                 �Yu@`��>�ϗ?/            @U@       �       �                 ��L@`���i��?             F@       ������������������������       �                     C@        �       �                    >@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �D@        �       �                 �|�=@�����?'            �R@       �       �                 pf� @ pƵHP�?             J@        ������������������������       �                     9@        �       �                   �;@ 7���B�?             ;@       �       �                 @3�!@$�q-�?             *@        �       �                   �7@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        �       �                 �y'"@���!pc�?             6@       �       �                 @3�@���N8�?             5@        �       �                   �?@�q�q�?             (@        ������������������������       �                     �?        �       �                   �A@���|���?             &@        ������������������������       �      �?             @        ������������������������       �����X�?             @        ������������������������       �                     "@        ������������������������       �                     �?        �       �                 ���#@�<ݚ�?             2@        ������������������������       �                      @        �       �                    3@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                   @C@D^��#��?1            �T@       �       �                    #@)O���?*             R@        �       �                    �?r�q��?             (@       �       �                    @����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��S���?#             N@        �       �                 ��$1@�㙢�c�?             7@       �       �                 ��.@�	j*D�?	             *@        �       �                    �?z�G�z�?             @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    @���"͏�?            �B@       �       �                    9@@�0�!��?             A@        ������������������������       �                     $@        �       �                   @@@      �?             8@       �       �                 �T)D@�q�q�?             2@       �       �                 ��2@d}h���?	             ,@       �       �                    �?      �?              @        ������������������������       �                     �?        �       �                 @3�/@և���X�?             @        ������������������������       �                     �?        �       �                 �|�;@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�;@      �?             @        ������������������������       �                      @        �       �                 �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    @ >�֕�?            �A@        ������������������������       �                     $@        �       �                    @HP�s��?             9@       �       �                 ��T?@�r����?             .@       ������������������������       �                     $@        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������.���|�?ӣ���?�z�G��?���(\��?�qa�?p�GOp�?�������?�������?����?����Ǐ�?      �?                      �?333333�?�������?      �?      �?]t�E]�?�E]t��?      �?        UUUUUU�?�������?333333�?ffffff�?      �?      �?      �?      �?      �?                      �?              �?      �?                      �?      �?        I�$I�$�?۶m۶m�?�,d!Y�?�Mozӛ�?��N��N�?�؉�؉�?q=
ףp�?{�G�z�?/�袋.�?F]t�E�?      �?      �?              �?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?333333�?�������?�������?�������?              �?      �?        wwwwww�?�?      �?        ]t�E]�?F]t�E�?�������?UUUUUU�?      �?              �?      �?              �?      �?        �������?333333�?              �?      �?        �������?�������?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        GX�i���?���=��?vb'vb'�?;�;��?+l$Za�?�'�K=�?      �?        ï�Dz��?z�rv��?۶m۶m�?%I�$I��?(�����?�k(���?              �?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?              �?�q�q�?�q�q�?�������?�������?      �?                      �?              �?      �?        �q�q�?�q�q�?              �?�������?�������?      �?      �?              �?      �?                      �?�؉�؉�?;�;��?)\���(�?���Q��?�������?UUUUUU�?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?                      �?      �?              �?              �?        {	�%���?������?              �?9��8���?�8��8��?              �?      �?        �����?6�&f�1�?}g���Q�?1���\�?B����?���+��?p�}��?Hp�}�?;�;��?�;�;�?L� &W�?m�w6�;�?�?�?              �?d!Y�B�?ӛ���7�?�������?333333�?              �?      �?                      �?ى�؉��?;�;��?              �?r�q��?�q�q�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?�������?              �?      �?              �?        z����?�/�ظ?��QNG9�?\cq��5�?      �?        �S� w��?�be�F�?              �?�n�Wc"�?���@��?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?��+j�?[�R�֯�?��o��o�?�A�A�?۶m۶m�?�$I�$I�?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?      �?/�袋.�?F]t�E�?xxxxxx�?�?      �?        �m۶m��?�$I�$I�?              �?ى�؉��?�؉�؉�?      �?              �?      �?      �?              �?        ���c�?��N�©?�������?�?F]t�E�?F]t�E�?      �?        �������?UUUUUU�?      �?                      �?      �?        �Ϻ���?v�)�Y7�?'vb'vb�?;�;��?      �?        	�%����?h/�����?�؉�؉�?;�;��?�������?UUUUUU�?      �?                      �?      �?              �?        F]t�E�?t�E]t�?�a�a�?��y��y�?�������?�������?              �?]t�E]�?F]t�E�?      �?      �?�m۶m��?�$I�$I�?      �?                      �?9��8���?�q�q�?      �?        333333�?�������?              �?      �?        ,Q��+�?�]�ڕ��?��8��8�?9��8���?UUUUUU�?�������?�$I�$I�?�m۶m��?              �?      �?                      �?�?�������?d!Y�B�?�7��Mo�?;�;��?vb'vb'�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?        �$I�$I�?�m۶m��?              �?      �?                      �?v�)�Y7�?*�Y7�"�?ZZZZZZ�?�������?      �?              �?      �?UUUUUU�?UUUUUU�?I�$I�$�?۶m۶m�?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?      �?                      �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?                      �?      �?        ��+��+�?�A�A�?      �?        q=
ףp�?{�G�z�?�������?�?      �?        333333�?�������?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJf��'hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       f                    �?>AU`�z�?�           8�@               _                 ��R@Ft����?�            �n@              
                    @�sD>�@�?�            �h@                                    @���7�?             6@        ������������������������       �                     ,@                                   @      �?              @       ������������������������       �                     @               	                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   (@�.�+��?t            �e@        ������������������������       �                      @               ^                    @rp��P��?o            �d@              =                 ��.@�G�z.�?l             d@                                    @�w�r��?4            @S@                                  �J@      �?             8@                               `f�)@���7�?             6@        ������������������������       �                     $@                                  �*@�8��8��?             (@                                  �?      �?              @                                 @<@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @               2                    �?X�Emq�?#            �J@              -                 �̌@�(�Tw��?            �C@              ,                    @�חF�P�?             ?@              !                   �3@��<b���?             7@                                 ��@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        "       '                 pff@r�q��?             2@        #       $                    �?���Q��?             @        ������������������������       �                     �?        %       &                 �|Y:@      �?             @       ������������������������       �                      @        ������������������������       �                      @        (       )                    �?$�q-�?             *@       ������������������������       �                     "@        *       +                   �7@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        .       /                 ��&@      �?              @        ������������������������       �                     @        0       1                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        3       4                 �!@؇���X�?             ,@        ������������������������       �                     �?        5       <                    �?$�q-�?             *@       6       ;                    �?ףp=
�?             $@       7       :                 ���,@      �?             @       8       9                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        >       ]                 ��qB@���O1��?8            �T@       ?       T                    �?     ��?+             P@       @       M                     @f1r��g�?"            �J@       A       F                    �?�L���?            �B@        B       E                     �?z�G�z�?             $@        C       D                 03�=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        G       L                    �? 7���B�?             ;@       H       I                   �E@��S�ۿ?             .@       ������������������������       �                     &@        J       K                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        N       O                    �?     ��?             0@        ������������������������       �                     @        P       Q                 �|�;@      �?             $@        ������������������������       �                     @        R       S                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        U       V                 ��97@���|���?	             &@        ������������������������       �                     @        W       X                     @      �?              @        ������������������������       �                      @        Y       Z                 X��@@�q�q�?             @        ������������������������       �                     @        [       \                   @C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     @        `       a                    �?@��8��?             H@       ������������������������       �                     D@        b       c                    �?      �?              @        ������������������������       �                     �?        d       e                    )@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        g       n                    @��QT(��?.           0}@        h       i                    @z�G�z�?             .@       ������������������������       �                     &@        j       m                    @      �?             @       k       l                 ���A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        o                         �R@p�̔B��?#           @|@       p       �                     �?P��sg��?"            |@        q       �                    �?     ��?@             X@        r       �                 p�w@H�z�G�?             D@       s       �                    �?؀�:M�?            �B@       t       �                 p"�X@П[;U��?             =@       u       �                    J@\X��t�?             7@       v       y                 ���<@     ��?
             0@        w       x                   @@@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        z                           �?$�q-�?             *@       {       |                 X�l@@�����H�?             "@        ������������������������       �                     @        }       ~                    C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �\@      �?              @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?����X�?*             L@        ������������������������       �                      @        �       �                   �<@l��
I��?)             K@        �       �                 `f�D@z�G�z�?             @       ������������������������       �                     @        �       �                    0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @@ \� ���?$            �H@        �       �                    K@\X��t�?             7@       �       �                 03:@      �?             4@        ������������������������       �                     @        �       �                    H@�θ�?
             *@       �       �                   @=@�q�q�?             "@       �       �                 �|�?@և���X�?             @        ������������������������       �                     �?        �       �                    D@�q�q�?             @        ������������������������       �                     @        �       �                 `f�;@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��9L@$�q-�?             :@       ������������������������       �                     2@        �       �                    G@      �?              @       �       �                 ��n^@���Q��?             @       �       �                 `f�N@�q�q�?             @        ������������������������       �                     �?        �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �                          �?p���87�?�             v@       �                          �?L��rH�?�            Pu@       �       �                     @�^����?�            pt@        �       �                   �*@�˹�m��?1             S@       �       �                    �?(L���?            �E@        ������������������������       �                     �?        �       �                 `fF)@؇���X�?             E@       �       �                    5@�C��2(�?             6@        �       �                   �2@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        �       �                 �|�<@z�G�z�?             4@        ������������������������       �                     $@        �       �                 �|�=@���Q��?             $@        ������������������������       �                      @        �       �                    @@      �?              @        ������������������������       �                      @        �       �                    C@�q�q�?             @        ������������������������       �                     �?        �       �                   �F@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                    �@@        �                       �T)D@ ���1��?�            `o@       �       �                 �?�@��� ��?�             o@       �       �                   �<@Du9iH��?U             `@        �       �                    �?�O4R���?!            �J@       �       �                   �4@���J��?             �I@        �       �                 P�@�X�<ݺ?
             2@        ������������������������       �                     $@        �       �                 �Y�@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �@@        ������������������������       �                      @        �       �                    �?�KM�]�?4             S@        �       �                 �|Y=@�8��8��?             8@        ������������������������       �                     �?        �       �                 �|�=@�nkK�?             7@       �       �                 ���@      �?             0@        ������������������������       �                     @        �       �                   @@�C��2(�?             &@       ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ���@ȵHPS!�?&             J@        ������������������������       �                     8@        �       �                    �?d}h���?             <@       �       �                 �Yu@�<ݚ�?             ;@       �       �                    B@ҳ�wY;�?             1@       �       �                   �?@և���X�?	             ,@       �       �                 �|Y=@�q�q�?             (@        ������������������������       �                     �?        �       �                    �?���!pc�?             &@       �       �                 ��(@      �?              @       ������������������������       �z�G�z�?             @        ������������������������       �                     @        �       �                 �|Y>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        �       �                 @3�@p�5�9��?K            �]@        �       �                   �?@�C��2(�?             &@        ������������������������       �                     @        �       �                   �A@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        �       
                   �?�e/
�?F             [@       �                       ��q1@W�!?�??            �X@       �                       �&�)@<����?<            �W@       �       �                   �3@�KM�]�?1             S@        �       �                 pf� @�q�q�?
             .@        �       �                   �1@�q�q�?             @        ������������������������       �      �?              @        ������������������������       �      �?             @        �       �                    ,@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���"@�.ߴ#�?'            �N@       ������������������������       �                     �J@                                 �<@      �?              @       ������������������������       �                     @                              �|Y=@      �?             @        ������������������������       �                      @                              �|�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@              	                   ;@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 �?�q�q�?             "@        ������������������������       �                     �?                                 +@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     *@        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?C��6�S�?�S\2��?T�r
^N�?և���X�?F]t�E�?�.�袋�?              �?      �?      �?              �?      �?      �?      �?                      �?�2)^ �?�f��o�?      �?        �7�:���?>�b���?ffffff�?ffffff�?
qV~B��?{����1�?      �?      �?F]t�E�?�.�袋�?              �?UUUUUU�?UUUUUU�?      �?      �?�������?�������?      �?                      �?              �?              �?      �?        �}�	��?5�x+��?� � �?�o��o��?��RJ)��?�Zk����?��Moz��?��,d!�?�������?333333�?              �?      �?        UUUUUU�?�������?�������?333333�?              �?      �?      �?              �?      �?        ;�;��?�؉�؉�?              �?      �?      �?              �?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?�������?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        ���ˊ��?P�M�_�?      �?      �?�x+�R�?�!5�x+�?L�Ϻ��?}���g�?�������?�������?      �?      �?      �?                      �?              �?h/�����?	�%����?�?�������?              �?      �?      �?              �?      �?                      �?      �?      �?              �?      �?      �?      �?        �$I�$I�?�m۶m��?              �?      �?        F]t�E�?]t�E]�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?�$I�$I�?۶m۶m�?      �?                      �?�p�RS��?M<洲�?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        X驅���?�ZX驅�?hE#߼�?b�r���?      �?      �?ffffff�?333333�?E>�S��?v�)�Y7�?�{a���?��=���?��Moz��?!Y�B�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?;�;��?�؉�؉�?�q�q�?�q�q�?              �?      �?      �?      �?                      �?              �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�m۶m��?�$I�$I�?      �?        Lh/����?h/�����?�������?�������?              �?      �?      �?              �?      �?        
^N��)�?և���X�?!Y�B�?��Moz��?      �?      �?      �?        �؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?        �؉�؉�?;�;��?      �?              �?      �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        T���5K�?a��S��?'�p�	'�?�{�Ǿ?οV���?� ����?��P^Cy�?^Cy�5�?⎸#��?w�qG��?      �?        ۶m۶m�?�$I�$I�?]t�E�?F]t�E�?333333�?�������?      �?                      �?      �?        �������?�������?      �?        333333�?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?              �?        �';r���?�`7>��?�{����?�B!��?qG�w��?w�qGܱ?:�&oe�?�x+�R�?______�?�?��8��8�?�q�q�?      �?              �?      �?              �?      �?              �?              �?        �k(���?(�����?UUUUUU�?UUUUUU�?              �?�Mozӛ�?d!Y�B�?      �?      �?      �?        ]t�E�?F]t�E�?�������?UUUUUU�?      �?              �?        ��N��N�?�؉�؉�?      �?        I�$I�$�?۶m۶m�?9��8���?�q�q�?�������?�������?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?F]t�E�?t�E]t�?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?              �?        �����?�O��O��?F]t�E�?]t�E�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?_B{	�%�?	�%��о?�v���?1ogH�۹?���%N�?�X�0Ҏ�?�k(���?(�����?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?      �?�q�q�?�q�q�?              �?      �?        �K�`m�?XG��).�?      �?              �?      �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?              �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJy"rhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                    �?�s�ˈ.�?�           8�@              �                    �?�(s�=�?a           �@                                   �?~6�����?           pz@                                  �9@�N��D�?<            �U@                                   �?�c�Α�?             =@        ������������������������       �                      @                                  �3@�ՙ/�?             5@                                hfF"@ףp=
�?             $@        	       
                 P��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                n"BT@���|���?	             &@                                 �7@�<ݚ�?             "@                               @3�@�q�q�?             @        ������������������������       �                     �?                                `fV$@z�G�z�?             @       ������������������������       �                     @                                  �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                �&�@��ϭ�*�?'             M@                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                  @B@ 7���B�?$             K@       ������������������������       �                    �D@                                `f�&@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        !       �                 ��q1@H��?"�?�             u@       "       #                 ���@���	���?�             q@        ������������������������       �                     =@        $       %                 ��@`U���H�?�            �n@        ������������������������       �                      @        &       5                    �?�Zl�i��?�            `n@        '       (                     @      �?             8@        ������������������������       �                     @        )       *                 ���@R���Q�?             4@        ������������������������       �                     @        +       ,                   �5@z�G�z�?             .@        ������������������������       �                     �?        -       2                   @@؇���X�?
             ,@       .       /                 �|=@ףp=
�?             $@        ������������������������       �                     @        0       1                 �|�=@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        3       4                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        6       �                   @F@����1�?�            `k@       7       J                     @     ��?~             h@        8       C                   �@@r�q��?             B@       9       <                    5@HP�s��?             9@        :       ;                   �2@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        =       >                   �'@���N8�?             5@        ������������������������       �                      @        ?       @                 �|�<@$�q-�?	             *@       ������������������������       �                     $@        A       B                 �|�=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        D       E                   @A@���|���?             &@        ������������������������       �      �?             @        F       G                   �'@����X�?             @        ������������������������       �                     �?        H       I                   @D@�q�q�?             @        ������������������������       �                      @        ������������������������       �      �?             @        K       T                    �?4��?�?h            �c@        L       M                 ���@�KM�]�?             3@        ������������������������       �                     @        N       S                 ��(@      �?             0@       O       P                 �|Y=@�r����?
             .@        ������������������������       �                     �?        Q       R                 X��A@@4և���?	             ,@       ������������������������       ��8��8��?             (@        ������������������������       �                      @        ������������������������       �                     �?        U       d                   �:@���	���?Z             a@        V       c                   �3@����˵�?'            �M@        W       b                 0S5 @؇���X�?             5@       X       _                   �2@���!pc�?
             &@       Y       \                    1@�q�q�?             @        Z       [                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ]       ^                 ��@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        `       a                 �?�@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     C@        e       �                   @@@�ݜ�?3            �S@       f       i                   �;@��.��?+            �N@        g       h                 �� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        j       y                 ��) @@�r-��?)            �M@       k       p                   �>@�C��2(�?             F@       l       o                 �?$@��?^�k�?            �A@        m       n                 pf�@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ?@        q       r                 �&B@�q�q�?             "@        ������������������������       �                     �?        s       t                   �?@      �?              @        ������������������������       �                     �?        u       v                   �@����X�?             @        ������������������������       �                     �?        w       x                 �?�@r�q��?             @        ������������������������       �                     �?        ������������������������       �z�G�z�?             @        z       {                   �<@�q�q�?
             .@        ������������������������       �                     @        |       �                    ?@      �?             $@       }       �                 ���(@      �?              @       ~       �                 ���"@����X�?             @              �                 �|Y=@      �?             @        ������������������������       �                     �?        �       �                 pf� @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     ;@        �       �                   �4@¦	^_�?)             O@        ������������������������       �                     @        �       �                   �R@0B��D�?(            �M@       �       �                   @J@�MWl��?'            �L@       �       �                    �?P����?             C@        �       �                 p�w@և���X�?             @       �       �                 ��tA@�q�q�?             @        �       �                 ���<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �>@�4�����?             ?@       �       �                 `fF:@X�<ݚ�?             2@        ������������������������       �                     @        �       �                   @=@և���X�?	             ,@       �       �                    H@X�<ݚ�?             "@       �       �                 �|�<@����X�?             @        ������������������������       �                     �?        �       �                 X��B@r�q��?             @        ������������������������       �                      @        �       �                 `f�;@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @>@z�G�z�?             @       �       �                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                      @8�Z$���?	             *@       �       �                   �B@�C��2(�?             &@        �       �                 �|�<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                      @        �       �                    �?�U���?I             _@        �       �                    �?�ՙ/�?             E@       �       �                   �-@�����H�?             2@        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�<@      �?             0@        ������������������������       �                     @        �       �                      @ףp=
�?	             $@        ������������������������       �                     @        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    G@�q�q�?             8@       �       �                    :@�q�q�?             5@        �       �                   �5@z�G�z�?             @        �       �                    .@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �7@     ��?             0@        �       �                    �?և���X�?             @        ������������������������       �                     @        �       �                    /@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �       �                    @������?+            �T@       �       �                    �?d�� z�?*            @T@        �       �                   �7@���Q��?            �A@        �       �                 ���.@�q�q�?	             5@        ������������������������       �                     @        �       �                     @     ��?             0@        ������������������������       �                     �?        �       �                 �|�;@��S���?             .@        ������������������������       �                     @        �       �                 �|Y>@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             ,@        �       �                 ��9L@�nkK�?             G@       ������������������������       �                     E@        �       �                     �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �8@      �?g            �d@        �       �                   �2@      �?3             T@       �       �                     @|��?���?%             K@        ������������������������       �        
             *@        �       �                     @��]�T��?            �D@        �       �                    @���|���?             6@       ������������������������       �                     *@        �       �                    #@�����H�?             "@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �0@�}�+r��?             3@       ������������������������       �                     2@        ������������������������       �                     �?        �       �                    �?8�Z$���?             :@       �       �                     @�����?
             5@       ������������������������       �                     1@        �       �                   �6@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                     @���Q��?             @       �       �                    �?�q�q�?             @       �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �                       @�:x@�ՙ/�?4             U@       �       �                 ��-@gO�~k�?3            @T@        ������������������������       �                     @                               ��.@X���[�?-            �R@                                 �?      �?              @        ������������������������       �                     @                              �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              	                    @��y�:�?)            �P@                                �?��c:�?             G@        ������������������������       �                     3@        ������������������������       �                     ;@        
                         �?؇���X�?             5@        ������������������������       �                     �?                                 @ףp=
�?             4@                                �?�IєX�?             1@                              ���5@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                @C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub��������������0Ȍ��?��o��?�� �+�?0�z���?2�����?��&@z��?�2)^ �?�~�u�7�?�{a���?5�rO#,�?              �?�a�a�?�<��<��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?]t�E]�?F]t�E�?9��8���?�q�q�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?              �?      �?              �?                      �?|a���?����=�?      �?      �?              �?      �?        h/�����?	�%����?              �?;�;��?;�;��?      �?                      �?�<��<��?1�0��?V��,���?P�9��J�?      �?        �[���?d �?�*�?              �?�"e����?�����H�?      �?      �?      �?        333333�?333333�?      �?        �������?�������?              �?۶m۶m�?�$I�$I�?�������?�������?      �?        �������?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?        �Ν;w��?Ĉ#F��?     ��?      �?�������?UUUUUU�?q=
ףp�?{�G�z�?      �?      �?      �?              �?      �?��y��y�?�a�a�?      �?        �؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?        ]t�E]�?F]t�E�?      �?      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?�N��N��?ى�؉��?�k(���?(�����?      �?              �?      �?�������?�?              �?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?        V��,���?P�9��J�?W'u_�?��/���?۶m۶m�?�$I�$I�?F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?                      �?      �?              �?        \��[���?�i�i�?�����?������?      �?      �?      �?                      �?'u_�?��c+���?]t�E�?F]t�E�?_�_��?�A�A�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?�$I�$I�?�m۶m��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?              �?              �?        ��Zk���?�RJ)���?              �?�A�I��?��}ylE�?:��,���?�YLg1�?�P^Cy�?Q^Cy��?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?���Zk��?��RJ)��?r�q��?�q�q�?      �?        ۶m۶m�?�$I�$I�?r�q��?�q�q�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?      �?      �?                      �?              �?;�;��?;�;��?]t�E�?F]t�E�?      �?      �?              �?      �?              �?              �?      �?      �?                      �?      �?                      �?c�1��?�9�s��?�a�a�?�<��<��?�q�q�?�q�q�?      �?      �?              �?      �?              �?      �?              �?�������?�������?              �?�������?�������?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?      �?      �?�$I�$I�?۶m۶m�?      �?              �?      �?      �?                      �?      �?                      �?�v%jW��?��+Q��?��"e���?x�5?,�?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        �?�������?      �?        333333�?ffffff�?              �?      �?                      �?�Mozӛ�?d!Y�B�?      �?              �?      �?              �?      �?                      �?      �?      �?      �?      �?	�%����?{	�%���?              �?KԮD�J�?jW�v%j�?F]t�E�?]t�E]�?              �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?        �5��P�?(�����?      �?                      �?;�;��?;�;��?�a�a�?=��<���?              �?      �?      �?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?�<��<��?�a�a�?�n���?��"e���?      �?        ��:m��?�X�%��?      �?      �?              �?      �?      �?              �?      �?        �@��~�?~5&��?-d!Y��?�7��Mo�?              �?      �?        ۶m۶m�?�$I�$I�?              �?�������?�������?�?�?�q�q�?�q�q�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�A�'hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       P                    �?>AU`�z�?�           8�@               G                    @ƆQ����?�            �n@              @                    �?:	��ʵ�?�             l@                                  �?��K�# �?z            �g@                                  �2@`2U0*��?0            �R@                                P��+@8�Z$���?	             *@        ������������������������       �                     @               	                     @�q�q�?             @        ������������������������       �                     @        
                          �-@�q�q�?             @        ������������������������       �                     �?                                  �0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 S�-@0�z��?�?'             O@                                �Q,@���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        ������������������������       �                     D@               ?                    �?�'�f7��?J             ]@              $                     @4�^o�]�?G            @\@              #                  �v7@�}�+r��?0             S@                                   �2@PN��T'�?             ;@                                 �*@�8��8��?             8@                               `f&'@�����?             5@                                  �J@      �?              @       ������������������������       �                     @        ������������������������       �                     �?                                   :@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @        !       "                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �H@        %       :                    �?��%��?            �B@       &       9                   @B@l��[B��?             =@       '       8                   �@@
j*D>�?             :@       (       3                    ;@
;&����?             7@       )       *                   �2@ҳ�wY;�?             1@        ������������������������       �                     �?        +       2                 pf� @     ��?             0@       ,       1                   �8@�8��8��?             (@       -       .                   �6@؇���X�?             @       ������������������������       �                     @        /       0                 @3�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        4       5                 �|Y>@r�q��?             @        ������������������������       �                     @        6       7                 ��*@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ;       <                    7@      �?              @        ������������������������       �                     @        =       >                    >@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        A       B                    @��.k���?             A@        ������������������������       �                     @        C       D                     @����"�?             =@       ������������������������       �        
             0@        E       F                    )@8�Z$���?	             *@        ������������������������       �                      @        ������������������������       �                     &@        H       K                    @�S����?             3@        I       J                 ��T?@      �?             @       ������������������������       �                      @        ������������������������       �                      @        L       M                    4@��S�ۿ?	             .@       ������������������������       �                     (@        N       O                 ���d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        Q       �                    �?�ۨ� ��?&           0}@        R                           �?�q�q�?1            @T@       S       x                    �?V������?.            �R@       T       e                     �?R=6�z�?&            @P@        U       d                    N@      �?             4@       V       c                    C@      �?             0@       W       ^                 �|�=@�eP*L��?             &@       X       Y                   �9@և���X�?             @        ������������������������       �                     �?        Z       [                 ��2>@�q�q�?             @        ������������������������       �                     @        \       ]                 �M@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        _       `                   @@@      �?             @        ������������������������       �                      @        a       b                 03�@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        f       u                 83�0@z�G�z�?            �F@       g       l                   �6@z�G�z�?             D@        h       i                    0@�q�q�?             @        ������������������������       �                      @        j       k                 ��y@      �?             @        ������������������������       �                      @        ������������������������       �                      @        m       t                 �|�=@l��\��?             A@       n       o                 �|=@R���Q�?             4@        ������������������������       �                     @        p       q                 ���@d}h���?             ,@        ������������������������       �                     @        r       s                 p&�@�z�G��?             $@       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     ,@        v       w                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        y       |                      @�q�q�?             "@       z       {                 �̾w@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        }       ~                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     �?����X�?             @        ������������������������       �                     �?        �       �                    *@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?$�D�B{�?�             x@        �       �                    @�C��2(�?            �@@       �       �                 �|Y=@ȵHPS!�?             :@        ������������������������       �                      @        �       �                    �? �q�q�?             8@       ������������������������       �                     7@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    #@�����?�            v@        �       �                    @r٣����?            �@@       ������������������������       �        	             7@        �       �                    @z�G�z�?             $@       ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?     ��?�             t@       �       �                    �?<��\�:�?�            �r@       �       �                 ��$:@�+�$f��?�            `r@       �       �                     �?�XinD��?�            �m@        ������������������������       �                     $@        �       �                 ���@�J��?�            �l@        ������������������������       �                     B@        �       �                   �>@h2��v�?}             h@       �       �                     @�}�+r��?V            �`@        ������������������������       �        
             .@        �       �                 ���@�1e�3��?L            �]@        ������������������������       �                      @        �       �                 �?$@���"�?K             ]@        �       �                    �?ףp=
�?             4@       �       �                 �|�;@�KM�]�?             3@       ������������������������       �                     &@        �       �                 ��,@      �?              @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                 @3�@      �??             X@        ������������������������       �                    �A@        �       �                    �?�.ߴ#�?'            �N@       �       �                 @�!@�}�+r��?%            �L@       �       �                 ��) @�C��2(�?            �@@       �       �                   �2@ �q�q�?             8@        �       �                    1@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �       �                 0SE @�<ݚ�?             "@        ������������������������       �                     �?        �       �                 pf� @      �?              @        ������������������������       �                     @        �       �                    8@z�G�z�?             @        ������������������������       �                     @        �       �                 �|Y<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        ������������������������       �                     @        �       �                 @3�@R���Q�?'             N@        �       �                 �?�@�����?
             3@       �       �                   �@�����H�?             "@       �       �                 �&B@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �?@      �?             $@        ������������������������       �                     @        �       �                   �A@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                   �'@��p\�?            �D@        ������������������������       �                     3@        �       �                   @A@��2(&�?             6@        �       �                    1@�q�q�?             @        ������������������������       �      �?             @        ������������������������       �                      @        �       �                   �*@      �?             0@        �       �                   �F@z�G�z�?             @        �       �                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                      @�2�o�U�?&            �K@       �       �                    �?      �?#             H@       �       �                   �;@�t����?             A@        ������������������������       �                     �?        �       �                   �>@���!pc�?            �@@       �       �                    K@�G�z��?             4@       �       �                   @>@�n_Y�K�?
             *@       �       �                 03k:@      �?             $@        ������������������������       �                      @        �       �                   `G@      �?              @       �       �                 X��B@r�q��?             @        ������������������������       �                      @        �       �                 `f�;@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    R@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        �       �                 03�U@؇���X�?	             ,@       �       �                   �E@$�q-�?             *@       �       �                  x#J@r�q��?             @        ������������������������       �                     @        �       �                 `�iJ@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    >@����X�?             @       �       �                    ;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���S@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     2@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������.���|�?ӣ���?�}�K�`�?�`mާ�?l�l��?��O��O�?kP<�q�?�밄���?{�G�z�?���Q��?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �B!��?|���{�?F]t�E�?�.�袋�?              �?      �?                      �?5�rO#,�?sO#,�4�?�|٠��?}٠ɗ�?(�����?�5��P�?h/�����?&���^B�?UUUUUU�?UUUUUU�?�a�a�?=��<���?      �?      �?              �?      �?        ;�;��?�؉�؉�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?}���g�?���L�?GX�i���?���=��?;�;��?b'vb'v�?�Mozӛ�?Y�B��?�������?�������?      �?              �?      �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?              �?333333�?�������?      �?                      �?              �?�?�������?      �?        �i��F�?	�=����?              �?;�;��?;�;��?              �?      �?        (������?^Cy�5�?      �?      �?      �?                      �?�������?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�P��=��?��9��?UUUUUU�?UUUUUU�?�g�`�|�?o0E>��?Wj�Vj��?S+�R+��?      �?      �?      �?      �?t�E]t�?]t�E�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?              �?      �?              �?      �?                      �?      �?        �������?�������?ffffff�?ffffff�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?------�?�������?333333�?333333�?      �?        I�$I�$�?۶m۶m�?      �?        ffffff�?333333�?      �?      �?      �?              �?        333333�?�������?              �?      �?        UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?        �����?�?�#%��?]t�E�?F]t�E�?��N��N�?�؉�؉�?              �?�������?UUUUUU�?      �?                      �?      �?        W�đ���?�����?|���?>���>�?              �?�������?�������?      �?        333333�?�������?      �?              �?      �?              �?      �?             ��?      �?b*1��J�?�vV;��?�Cc}h�?/�����?�Y���?30]�X#�?      �?        �����?t�?;��?      �?        ~���X�?��H	9�?�5��P�?(�����?      �?        �/���?W'u_�?              �?X�i���?|a���?�������?�������?�k(���?(�����?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?        �K�`m�?XG��).�?�5��P�?(�����?]t�E�?F]t�E�?�������?UUUUUU�?      �?      �?      �?                      �?      �?        9��8���?�q�q�?              �?      �?      �?      �?        �������?�������?      �?              �?      �?              �?      �?              �?              �?        333333�?333333�?Q^Cy��?^Cy�5�?�q�q�?�q�q�?      �?      �?      �?                      �?      �?              �?      �?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?�]�ڕ��?��+Q��?      �?        ��.���?t�E]t�?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?�������?�������?      �?      �?      �?                      �?      �?              �?        ־a��?�S�<%��?      �?      �?�������?�������?              �?F]t�E�?t�E]t�?�������?�������?ى�؉��?;�;��?      �?      �?              �?      �?      �?�������?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?                      �?      �?        ۶m۶m�?�$I�$I�?�؉�؉�?;�;��?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������                           @�����?�           8�@               	                 03�=@���N8�?             E@                                  �?�nkK�?             7@                               ��*4@�IєX�?             1@       ������������������������       �        	             (@                                ���7@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        
                            @�\��N��?
             3@                                   �?      �?              @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                   �?���!pc�?             &@                                ��T?@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                   @؇���X�?             @                                  @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @               x                     @z/����?�           �@               o                   @N@4��@���?�            �r@              4                    �?ħ�,{��?�            �q@               )                   �B@����p�?Q             a@                                  �?x��B�R�?8            �V@        ������������������������       �                     <@               (                    �?���N8�?&            �O@               !                    �?��p\�?            �D@       ������������������������       �                     8@        "       #                     �?@�0�!��?
             1@        ������������������������       �                     @        $       '                   �;@      �?             (@        %       &                    7@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     6@        *       3                 ��A@���V��?            �F@        +       ,                    �?�q�q�?
             5@        ������������������������       �                     @        -       0                   �6@@�0�!��?	             1@       .       /                   �C@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        1       2                     �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     8@        5       Z                     �?V��~��?g            �b@       6       Q                    �?&:~�Q�?4             S@       7       F                  �>@0�� ��?+            �O@       8       9                 ��<:@l��[B��?             =@        ������������������������       �                      @        :       E                    K@����X�?             5@       ;       D                 ��=@r�q��?             2@       <       C                   `G@�q�q�?             "@       =       @                    �?      �?             @        >       ?                 ��";@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        A       B                   �C@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        G       H                   �7@�t����?             A@        ������������������������       �                      @        I       P                    �?      �?             @@       J       M                 �|�<@�8��8��?             8@        K       L                    :@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        N       O                 p�w@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                      @        R       Y                 Ј�U@�n_Y�K�?	             *@       S       X                   �E@      �?              @        T       W                   @B@      �?             @       U       V                   @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        [       n                    �?@-�_ .�?3            �R@       \       m                   �*@ 	��p�?'             M@       ]       d                   �@@�����?             E@       ^       c                    5@ ��WV�?             :@        _       `                   �2@      �?              @       ������������������������       �                     @        a       b                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        e       f                   �)@     ��?             0@        ������������������������       �                      @        g       l                   �F@      �?              @       h       k                   @D@      �?             @       i       j                   �A@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             0@        ������������������������       �                     0@        p       q                    �?؇���X�?             ,@        ������������������������       �                     @        r       w                     @"pc�
�?
             &@       s       t                    �?�<ݚ�?	             "@        ������������������������       �                     �?        u       v                   �R@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        y       �                    �?�zц��?�            w@        z       �                    �?)b���?F            �Z@       {       �                    �?҄��?.            �P@        |       }                 03�)@�g�y��?             ?@       ������������������������       �                     7@        ~                           �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?<=�,S��?            �A@       �       �                    ;@�\��N��?             3@       �       �                   �3@���|���?	             &@        ������������������������       �                     �?        �       �                 @q"@�z�G��?             $@       �       �                    8@�<ݚ�?             "@       ������������������������       �                     @        �       �                 �&B@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��� @      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �|�;@      �?             0@       �       �                   �3@�C��2(�?             &@        �       �                 �y�)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                     @���Q��?             @       �       �                 X�,C@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?� ��1�?            �D@        �       �                    +@�q�q�?             5@        ������������������������       �                     @        �       �                    7@��S���?	             .@        �       �                 ��'@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y=@�q�q�?             "@        ������������������������       �                     @        �       �                 �A7@      �?             @       �       �                 hV}1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 @34@P���Q�?             4@        �       �                 �|�:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        �       �                    #@��E���?�            `p@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                     @���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    @     p�?�             p@       �       �                    �?HP�s��?�            @o@       �       �                   @@@���X=P�?�            �n@       �       �                    �?��(!i�?y            �h@       �       �                 �?�@��0��?i            �e@       �       �                    �?@4և���?B             \@        �       �                 ���@����X�?             ,@        �       �                 �|�9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @8@���!pc�?             &@        ������������������������       �                      @        �       �                 �|=@�����H�?             "@        ������������������������       �                      @        �       �                 �|�=@؇���X�?             @       ������������������������       �r�q��?             @        ������������������������       �                     �?        �       �                    �?@9G��?:            �X@        �       �                  ��@�nkK�?             7@        ������������������������       �                     $@        �       �                 ��(@$�q-�?             *@       ������������������������       ��8��8��?             (@        ������������������������       �                     �?        �       �                   �@`2U0*��?.            �R@       �       �                   �?@��<D�m�?            �H@       �       �                 �|�<@`Ql�R�?            �G@       ������������������������       �                     C@        �       �                 �|Y>@�����H�?             "@       �       �                 pf�@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     :@        �       �                    �?R���Q�?'             N@        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 0SE @Ԫ2��?$            �L@       �       �                   �2@������?             >@        �       �                    1@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        �       �                 �|Y=@�<ݚ�?             ;@        ������������������������       �                     @        �       �                 ��) @�z�G��?             4@       �       �                 �|Y>@@�0�!��?
             1@       ������������������������       �                     $@        �       �                   �?@և���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     ;@        �       �                    �?�8��8��?             8@       �       �                    6@�t����?             1@        �       �                    3@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                    �H@        �       �                  �v6@z�G�z�?             @       ������������������������       �                     @        �       �                 �|�:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub������������������?��܍��?��y��y�?�a�a�?d!Y�B�?�Mozӛ�?�?�?              �?�������?�������?      �?                      �?              �?�5��P�?y�5���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?t�E]t�?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?        ,�����?��u<J�?�G�z�?�(\����?T�ik���?V0K���?�����Ҳ?�������?��?�����?              �?�a�a�?��y��y�?��+Q��?�]�ڕ��?              �?�������?ZZZZZZ�?              �?      �?      �?333333�?�������?              �?      �?                      �?              �?�>�>��?[�[��?UUUUUU�?UUUUUU�?      �?        �������?ZZZZZZ�?UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?              �?      �?                      �?c�/��b�?t�@�t�?�k(���?�k(����?�eY�eY�?�4M�4M�?GX�i���?���=��?      �?        �$I�$I�?�m۶m��?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?                      �?              �?      �?        <<<<<<�?�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?ffffff�?�������?      �?                      �?      �?        ى�؉��?;�;��?      �?      �?      �?      �?      �?      �?      �?                      �?              �?      �?                      �?S�n0E�?к����?������?�{a���?=��<���?�a�a�?O��N���?;�;��?      �?      �?      �?              �?      �?              �?      �?              �?              �?      �?      �?              �?      �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?              �?              �?        ۶m۶m�?�$I�$I�?      �?        /�袋.�?F]t�E�?9��8���?�q�q�?              �?      �?      �?      �?                      �?      �?        @��(��?o`E\��?����f��?��4>2��?N6�d�M�?�d�M6��?�B!��?��{���?              �?      �?      �?      �?                      �?�A�A�?X|�W|��?y�5���?�5��P�?F]t�E�?]t�E]�?      �?        333333�?ffffff�?�q�q�?9��8���?              �?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?      �?      �?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?333333�?      �?      �?              �?      �?                      �?������?������?UUUUUU�?UUUUUU�?      �?        �?�������?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?      �?                      �?      �?        ffffff�?�������?      �?      �?              �?      �?              �?        T���0�?�_�	)y�?      �?      �?      �?        �������?333333�?      �?              �?      �?              �?      �?             ��?      �?q=
ףp�?{�G�z�?�j򸳄�?]�l8bڳ?9/����?4և��и?6eMYS��?S֔5eM�?n۶m۶�?�$I�$I�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?        ������?9/���?�Mozӛ�?d!Y�B�?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?        ���Q��?{�G�z�?��S�r
�?և���X�?}g���Q�?W�+�ɕ?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?      �?                      �?      �?        333333�?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        $���>��?p�}��?wwwwww�?�?UUUUUU�?UUUUUU�?      �?      �?              �?9��8���?�q�q�?      �?        ffffff�?333333�?ZZZZZZ�?�������?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?<<<<<<�?�?333333�?�������?      �?                      �?      �?              �?              �?        �������?�������?      �?              �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJJ��hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM)hjh))��}�(h,h/h0M)��h2h3h4hph<�h=Kub������       �                     @�,�٧��?�           8�@                                   �?Y(���?�            �s@                                  �E@Du9iH��?L             `@                                   �?�f�¦ζ??            �Z@        ������������������������       �                     J@                                  �6@�C��2(�?!            �K@                                  �?��hJ,�?             A@              	                    �?д>��C�?             =@        ������������������������       �                     @        
                           <@���B���?             :@                                  �6@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @                                  �'@�IєX�?             1@        ������������������������       �                     @                                   1@$�q-�?             *@                                 �B@�C��2(�?             &@       ������������������������       �                     "@                                   D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@                                   �?"pc�
�?             6@                                83F@����X�?             @        ������������������������       �                      @        ������������������������       �                     @                                  @F@�r����?	             .@        ������������������������       �                      @        ������������������������       �                     *@                c                    �?�7����?s            �g@       !       "                   �1@4�2%ޑ�?X            �a@        ������������������������       �                     @        #       J                     �?H�V�e��?U             a@       $       I                    �?��Q���?0             T@       %       D                    �?�(�Tw��?/            �S@       &       ?                  �>@j�'�=z�?)            �P@       '       4                    D@��.k���?             A@       (       )                 ��I/@�q�q�?             5@        ������������������������       �                     @        *       +                    <@      �?
             0@        ������������������������       �                     @        ,       -                 �|Y=@z�G�z�?             $@        ������������������������       �                     �?        .       3                    �?�����H�?             "@        /       2                 X�,@@      �?             @       0       1                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        5       >                    R@8�Z$���?	             *@       6       =                   �J@�8��8��?             (@        7       8                 ��:@r�q��?             @        ������������������������       �                      @        9       <                 `f�;@      �?             @       :       ;                   @G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        @       C                 �|Y<@      �?             @@        A       B                   �9@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     <@        E       H                    �?�q�q�?             (@       F       G                   @B@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        K       L                    �? �Cc}�?%             L@        ������������������������       �                     @        M       `                   @D@���C��?"            �J@       N       _                   �3@�8��8��?             H@       O       P                    @������?            �D@        ������������������������       �                     @        Q       V                    5@�����H�?             B@        R       S                   �2@"pc�
�?             &@        ������������������������       �                     @        T       U                   �'@      �?              @       ������������������������       ����Q��?             @        ������������������������       �                     @        W       \                   �@@HP�s��?             9@       X       [                 �|�=@P���Q�?             4@       Y       Z                 �|Y=@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     $@        ]       ^                   @B@z�G�z�?             @       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        a       b                   @F@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        d       }                    �?�q�q�?             H@       e       l                    �?���Q��?            �F@        f       g                   �5@���|���?             &@        ������������������������       �                     @        h       i                 м{G@      �?              @        ������������������������       �                      @        j       k                 p"�X@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        m       z                     �?j���� �?             A@       n       u                 03�M@8�A�0��?
             6@        o       p                  x#J@���Q��?             $@        ������������������������       �                     @        q       r                    A@؇���X�?             @        ������������������������       �                     @        s       t                   �C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        v       w                    �?      �?             (@       ������������������������       �                     @        x       y                �G�:@@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        {       |                    :@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                     @        ~                           �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �0@L K6R�?	           �x@        �       �                   �-@~h����?(             L@       �       �                 @3�4@�q�����?#             I@        �       �                    @�+$�jP�?             ;@       ������������������������       �        	             (@        �       �                    �?�q�q�?             .@        �       �                 �&�)@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    $@�����H�?             "@        ������������������������       �                     @        �       �                 �y.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?���}<S�?             7@        ������������������������       �                     "@        �       �                    @؇���X�?             ,@        ������������������������       �                     @        �       �                    �?z�G�z�?	             $@       �       �                    @z�G�z�?             @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @z�G�z�?             @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �      �?              @        �       �                    �?�θ�?�             u@        �       �                 ��,#@fK!���?9            �V@        �       �                    �?6YE�t�?            �@@       �       �                  ��@r�q��?             >@       �       �                  s@؇���X�?             <@        ������������������������       �                     @        �       �                    �?"pc�
�?             6@       ������������������������       �        	             *@        �       �                 �&B@X�<ݚ�?             "@       �       �                 ���@      �?              @        �       �                 �|Y:@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    7@T����1�?#             M@        �       �                    �?$�q-�?             *@        �       �                  �#@      �?             @        ������������������������       �                      @        �       �                 �[$@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    @���Q��?            �F@       �       �                 ��.@�\��N��?             C@        �       �                    �?z�G�z�?             $@        ������������������������       �                     @        �       �                   �*@���Q��?             @       �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��Y7@և���X�?             <@       �       �                 �|�;@z�G�z�?	             .@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�	j*D�?             *@        ������������������������       �                     @        �       �                    @ףp=
�?             $@        ������������������������       �                     @        �       �                   @C@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �                         @@@l�ْ��?�            �n@       �                          �?8�Z$���?�            `h@       �                          �?�&U��y�?y            �f@       �       �                    �?t�6Z���?m            �d@        �       �                 ���@z�G�z�?            �A@        �       �                   �7@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 ��(@      �?             8@       �       �                 �Y�@�z�G��?             4@       �       �                    �?�<ݚ�?             "@       �       �                   �5@����X�?             @        ������������������������       �                     �?        �       �                 �|�:@r�q��?             @        ������������������������       �                      @        �       �                 �|�=@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|Y=@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �                         �?@��POc�?V            @`@       �       �                   �2@\#r��?P            �^@        �       �                 pf� @և���X�?             @        �       �                 ���@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �9@ج��w�?L            �\@        ������������������������       �        $             K@        �       �                 ��) @f>�cQ�?(            �N@       �       �                 �&B@ ���J��?            �C@        �       �                 �|�;@ףp=
�?             $@        ������������������������       �                      @        �       �                 �|Y>@      �?              @       �       �                 pf�@r�q��?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     =@        �                        pf� @���|���?             6@        ������������������������       �                      @                                �;@�z�G��?             4@        ������������������������       �                     @              
                �|Y=@      �?
             0@             	                ���)@�<ݚ�?             "@                              ���"@      �?             @        ������������������������       �                     �?                                �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                              P�@      �?              @        ������������������������       �                     @                              d�6@@���Q��?             @                             ��I @      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?                              �̌3@      �?             0@       ������������������������       �        	             (@                                 �?      �?             @                             03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                 �?X�Cc�?             ,@                              ��y&@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                  �? pƵHP�?'             J@        ������������������������       �                     "@        !      (                   �? qP��B�?            �E@       "      '                  �C@������?             B@        #      $                �?�@�}�+r��?             3@       ������������������������       �                     "@        %      &                @3�@ףp=
�?             $@        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M)KK��h2h3h4hVh<�h=Kub�������������&��jq�?:�g *�?��8BF�?�)���\�?w�qGܱ?qG�w��?�Ե��?��4>2��?              �?F]t�E�?]t�E�?�������?KKKKKK�?|a���?a���{�?              �?ى�؉��?��؉���?�q�q�?r�q��?              �?      �?        �?�?              �?;�;��?�؉�؉�?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?              �?              �?              �?F]t�E�?/�袋.�?�$I�$I�?�m۶m��?      �?                      �?�?�������?      �?                      �?]AL� &�?G}g����?�������?�A�A�?              �?iiiiii�?ZZZZZZ�?333333�?�������?�o��o��?� � �?�|���?|��|�?�������?�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?�������?�������?      �?        �q�q�?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?;�;��?;�;��?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?                      �?      �?              �?                      �?      �?      �?      �?      �?      �?                      �?      �?        �������?�������?�q�q�?r�q��?              �?      �?              �?              �?        %I�$I��?۶m۶m�?      �?        \�琚`�?"5�x+��?UUUUUU�?UUUUUU�?�|����?������?      �?        �q�q�?�q�q�?/�袋.�?F]t�E�?      �?              �?      �?333333�?�������?      �?        q=
ףp�?{�G�z�?ffffff�?�������?�������?�������?      �?                      �?      �?        �������?�������?      �?      �?      �?              �?        333333�?�������?              �?      �?        �������?�������?333333�?�������?]t�E]�?F]t�E�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?ZZZZZZ�?颋.���?/�袋.�?�������?333333�?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?      �?      �?        �������?333333�?              �?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�?��DO�?���@va�?�m۶m��?%I�$I��?�p=
ף�?���Q��?B{	�%��?/�����?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?        ӛ���7�?d!Y�B�?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?�������?�������?      �?      �?      �?                      �?      �?        �������?�������?      �?      �?              �?      �?              �?        UUUUUU�?�������?              �?      �?      �?ى�؉��?�؉�؉�?�����?q�p��?e�M6�d�?'�l��&�?UUUUUU�?�������?�$I�$I�?۶m۶m�?              �?F]t�E�?/�袋.�?              �?�q�q�?r�q��?      �?      �?�������?333333�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?              �?�FX�i��?�rO#,��?�؉�؉�?;�;��?      �?      �?      �?              �?      �?              �?      �?              �?        333333�?�������?y�5���?�5��P�?�������?�������?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ۶m۶m�?�$I�$I�?�������?�������?      �?      �?              �?      �?                      �?vb'vb'�?;�;��?              �?�������?�������?      �?        �������?UUUUUU�?              �?      �?              �?        ��1����?	9?��?;�;��?;�;��?�����?�1�����?X���oX�?��)A��?�������?�������?]t�E�?F]t�E�?              �?      �?              �?      �?ffffff�?333333�?9��8���?�q�q�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        ]t�E]�?F]t�E�?              �?      �?              �?        �����?�����?��:��?XG��).�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?        �%��~�?A�V���?      �?        ��!XG�?�u�y���?��-��-�?�A�A�?�������?�������?      �?              �?      �?�������?UUUUUU�?      �?              �?      �?      �?              �?        ]t�E]�?F]t�E�?              �?ffffff�?333333�?              �?      �?      �?9��8���?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?              �?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?              �?      �?      �?      �?              �?      �?              �?        %I�$I��?�m۶m��?�$I�$I�?�m۶m��?      �?                      �?      �?        'vb'vb�?;�;��?      �?        ��}A�?�}A_З?�q�q�?�q�q�?�5��P�?(�����?      �?        �������?�������?      �?      �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�U�uhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������       j                     @��t���?�           8�@                                   �?
֙g0��?�            �u@                                03�<@=0�_�?]             c@                                  �?$��$�L�?/            �S@                                   �?f1r��g�?!            �J@                                0#R;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        	                           �?�:pΈ��?             I@       
                           L@�X�<ݺ?             B@                                 �9@��?^�k�?            �A@                                   �?r�q��?             @        ������������������������       �                      @                                  �'@      �?             @        ������������������������       �                      @                                  �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     =@        ������������������������       �                     �?                                  �;@X�Cc�?             ,@                                  �9@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @                                   9@      �?              @        ������������������������       �                      @                                  �E@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     :@        ������������������������       �        .            �R@                9                 ��$:@�%����?u             h@        !       "                    #@ܷ��?��?6            �U@        ������������������������       �                     @        #       $                    �? 7���B�?3            @T@        ������������������������       �                     @        %       8                   �*@`2U0*��?/            �R@       &       3                   �D@��S�ۿ?            �F@       '       2                 �|�=@�}�+r��?             C@       (       -                 �|�<@�>����?             ;@       )       ,                    5@���N8�?             5@       *       +                    &@�8��8��?             (@        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     "@        .       /                     �?r�q��?             @        ������������������������       �                     �?        0       1                    @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             &@        4       5                 `f�)@؇���X�?             @        ������������������������       �                     �?        6       7                    G@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     >@        :       i                    @H(���o�??            �Z@       ;       f                    �?����3��?>             Z@       <       I                   �<@�X���?7             V@        =       B                   �8@�����?             3@        >       ?                    6@r�q��?             @        ������������������������       �                     @        @       A                 ���Q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        C       D                 `f�D@$�q-�?	             *@        ������������������������       �                     @        E       H                    �?r�q��?             @        F       G                 ��N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        J       K                 03k:@�G�5��?)            @Q@        ������������������������       �                      @        L       e                   �R@��ga�=�?(            �P@       M       d                    �?z�G�z�?'            @P@       N       [                  x;K@����|e�?!             K@       O       Z                  �>@�ݜ�?            �C@       P       Y                    �?���N8�?             5@       Q       X                   @>@�d�����?             3@       R       W                 `f�;@@�0�!��?
             1@       S       V                   �J@���!pc�?             &@        T       U                 X��B@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             2@        \       ]                 03�M@��S���?
             .@        ������������������������       �                     @        ^       _                    �?�<ݚ�?             "@        ������������������������       �                      @        `       c                    �?����X�?             @       a       b                   �G@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        g       h                    5@      �?             0@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        k       �                   @@@�|��gN�?�            �v@       l       �                    @      �?�            �r@       m       �                    �?��5Е��?�            �p@       n       q                 �ٝ@���?�            �l@        o       p                    �?@4և���?             E@        ������������������������       �                     @        ������������������������       �                    �C@        r       �                 ��@&�
�M�?}            �g@        s       z                  ��@X��ʑ��?            �E@        t       y                    �?b�2�tk�?
             2@       u       v                 �|Y:@�<ݚ�?             "@       ������������������������       �                     @        w       x                 @3�@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        {       |                    1@� �	��?             9@        ������������������������       �                     @        }       �                    �?      �?             6@       ~                        �|Y=@�G�z��?             4@        ������������������������       �                     @        �       �                    �?��.k���?             1@        ������������������������       �                     @        �       �                    �?ףp=
�?             $@       ������������������������       ������H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?V�a�� �?c             b@        �       �                    �?�n_Y�K�?             :@        �       �                 �|Y6@      �?              @        ������������������������       �                     @        �       �                    �?      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �:@r�q��?             2@        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|Y<@��S�ۿ?
             .@        ������������������������       �                     �?        �       �                    �?@4և���?	             ,@        ������������������������       �                     @        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��u}���?Q            �]@        �       �                    �?�eP*L��?             6@       �       �                    �?�G��l��?             5@       �       �                  sW@և���X�?	             ,@        ������������������������       �                      @        �       �                    =@�q�q�?             (@       �       �                    3@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �!@և���X�?             @        ������������������������       �                      @        �       �                 ���)@���Q��?             @        ������������������������       �                      @        �       �                 �|�7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��C@�^'�ë�?C            @X@       �       �                    �?���}<S�?A             W@       �       �                 �?�@�:�^���?@            �V@        ������������������������       �                     <@        �       �                 @3�@��� ��?,             O@        �       �                   �4@���Q��?             @        ������������������������       �                     �?        �       �                    :@      �?             @        ������������������������       �                     �?        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        �       �                 ���#@x�}b~|�?'            �L@       �       �                 ���"@X�EQ]N�?            �E@       �       �                 ��Y @ >�֕�?            �A@       �       �                   �2@�8��8��?             8@        �       �                    1@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     &@        �       �                    =@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             ,@        ������������������������       �                      @        �       �                    ;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�\��N��?             C@       �       �                    @ҳ�wY;�?             1@        ������������������������       �                     @        �       �                    �?�eP*L��?             &@       �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                 ��y&@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��\6@և���X�?
             5@       �       �                 �|Y=@���Q��?             .@       �       �                    9@ףp=
�?             $@       ������������������������       �                     @        �       �                  �1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?             @@        ������������������������       �                     (@        �       �                    @P���Q�?             4@        �       �                    �?      �?              @        ������������������������       �                     @        �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             (@        �       �                 @3�@��ɉ�?&            @P@        �       �                    �?��S�ۿ?             >@        ������������������������       �                     "@        �       �                 �?�@�����?             5@       ������������������������       �                     1@        ������������������������       �      �?             @        ������������������������       �                    �A@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������nԾ���?5"W��6�?ۜ��L|�?�������?p�pŪ?��S��S�?�3���?��]-n��?�x+�R�?�!5�x+�?UUUUUU�?UUUUUU�?              �?      �?        �Q����?��Q���?�q�q�?��8��8�?�A�A�?_�_��?UUUUUU�?�������?              �?      �?      �?              �?      �?      �?              �?      �?                      �?      �?        �m۶m��?%I�$I��?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?UUUUUU�?�������?              �?      �?                      �?              �?(b6�5�?aw&��+�?��=���?a���{�?              �?	�%����?h/�����?      �?        ���Q��?{�G�z�?�������?�?�5��P�?(�����?�Kh/��?h/�����?��y��y�?�a�a�?UUUUUU�?UUUUUU�?      �?      �?      �?              �?        �������?UUUUUU�?      �?        �������?�������?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        M0��>��?e�Cj���?��N��N�?'vb'vb�?]t�E�?�E]t��?^Cy�5�?Q^Cy��?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ;�;��?�؉�؉�?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?��v`��?�%~F��?              �?��[���?�1���?�������?�������?����K�?	�%����?\��[���?�i�i�?�a�a�?��y��y�?Cy�5��?y�5���?ZZZZZZ�?�������?F]t�E�?t�E]t�?�������?333333�?      �?                      �?      �?              �?                      �?      �?              �?        �������?�?              �?9��8���?�q�q�?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?      �?      �?              �?      �?              �?        ����?�?���� �?      �?      �?�jL�*�?*g���?�q�.�|�?�9E[�?n۶m۶�?�$I�$I�?              �?      �?        }g���Q�?1���\�?�}A_�?��}A�?�8��8��?9��8���?�q�q�?9��8���?              �?      �?      �?      �?                      �?      �?        )\���(�?�Q����?              �?      �?      �?�������?�������?              �?�������?�?              �?�������?�������?�q�q�?�q�q�?      �?              �?        ��{a�?a���{�?;�;��?ى�؉��?      �?      �?              �?      �?      �?      �?      �?      �?                      �?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?�������?�?      �?        n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?{1�z1��?:�:��?t�E]t�?]t�E�?1�0��?��y��y�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?      �?                      �?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        =�L�v��?���Id�?ӛ���7�?d!Y�B�?}�'}�'�?l�l��?      �?        �{����?�B!��?�������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?�YLg1�?Lg1��t�?w�qG�?qG�wĽ?��+��+�?�A�A�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?      �?                      �?      �?              �?        333333�?�������?              �?      �?        �5��P�?y�5���?�������?�������?              �?t�E]t�?]t�E�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�������?�������?              �?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?�������?333333�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?      �?      �?        ffffff�?�������?      �?      �?      �?        �������?�������?      �?              �?      �?      �?                      �?      �?        ?�?��? �����?�������?�?      �?        =��<���?�a�a�?      �?              �?      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW��]hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       B                    �?e�L��?�           8�@               =                    @��}� �?�            �o@              <                    @�9�K(��?�            �m@                                  �?��&y�X�?�             m@                                0Cd=@�C��2(�?8             V@                                 �B@��s����?             E@                                  �?�ݜ�?            �C@               	                   P,@����X�?             ,@        ������������������������       �                     @        
                        `�@1@      �?              @       ������������������������       �                     @        ������������������������       �                     @                                ���@`2U0*��?             9@        ������������������������       �                     �?        ������������������������       �                     8@        ������������������������       �                     @        ������������������������       �                     G@               !                   �9@~X�<��?Y             b@                                   �?�ՙ/�?&            �O@                                  �3@j���� �?             A@                                 �3@�q�q�?             >@        ������������������������       �                      @                                  �6@�C��2(�?             6@                                P @r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     $@        ������������������������       �                     @                                    @\-��p�?             =@       ������������������������       �                     3@                                 `f7@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        "       1                     @^�pӵL�?3            @T@       #       &                   �;@6uH���?&             O@        $       %                   �/@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        '       (                     �? ,��-�?$            �M@        ������������������������       �                     :@        )       0                   �*@<���D�?            �@@        *       -                 `f�)@����X�?             ,@       +       ,                   �J@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        .       /                   �A@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     3@        2       7                    �?�\��N��?             3@       3       6                    A@      �?              @       4       5                 �?�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        8       ;                 03�1@�eP*L��?             &@        9       :                   �D@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        >       ?                    0@      �?	             0@       ������������������������       �                     $@        @       A                      @�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        C       t                    �?��/T8�?"           �|@        D       I                   �2@¦	^_�?8            @W@        E       H                 pV�;@r�q��?             @        F       G                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        J       s                   �H@�6tT�.�?4            �U@       K       ^                     �?��It��?.            �S@        L       Y                  �	U@��
ц��?             :@       M       X                    �?�q�q�?
             .@       N       W                 X�l@@����X�?	             ,@       O       P                    9@���Q��?             $@        ������������������������       �                     @        Q       R                 �ܵ<@և���X�?             @        ������������������������       �                     �?        S       T                 �|Y<@�q�q�?             @        ������������������������       �                      @        U       V                 ��2>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        Z       [                 Ȫ�c@"pc�
�?             &@        ������������������������       �                     @        \       ]                 p�w@      �?             @        ������������������������       �                      @        ������������������������       �                      @        _       b                   �5@f1r��g�?             �J@        `       a                 �{@      �?             @        ������������������������       �                      @        ������������������������       �                      @        c       d                     @�q��/��?            �H@        ������������������������       �                     (@        e       r                    �?�MI8d�?            �B@       f       q                    �?l��\��?             A@       g       p                 @3s+@��a�n`�?             ?@       h       o                 �|�=@��S�ۿ?             >@       i       j                 ���@�����H�?             2@        ������������������������       �                     "@        k       l                 �|=@�<ݚ�?             "@        ������������������������       �                      @        m       n                   @@����X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        u       �                     �? M)���?�            �v@        v       �                 `��S@r�z-��?'            �J@       w       �                  i?@p�v>��?"            �G@        x       �                   @=@r�q��?             8@       y       �                   �K@d}h���?             ,@       z       {                 ��:@�z�G��?
             $@        ������������������������       �                     @        |       �                   `G@���Q��?             @       }       �                 `f�;@�q�q�?             @       ~                        �|�?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|Y=@z�G�z�?             $@        �       �                    <@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�LQ�1	�?             7@       ������������������������       �        	             &@        �       �                    F@      �?             (@       �       �                  x#J@      �?              @        ������������������������       �                      @        �       �                   �C@      �?             @       �       �                 `f�K@      �?             @        ������������������������       �                      @        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �T�I@��7H�?�            ps@       �       �                 �?�@؅�q(�?�            �r@        �       �                    �?T��,��?B            @Y@       �       �                    �?` A�c̭?A             Y@        �       �                 �|Y;@�nkK�?             7@        ������������������������       �                     �?        �       �                 �Y�@���7�?             6@        ������������������������       �                     @        �       �                    �?      �?	             0@       �       �                 ��(@��S�ۿ?             .@       ������������������������       �$�q-�?             *@        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�g<a�?4            @S@       �       �                 �|�<@�?�|�?2            �R@        ������������������������       �                     ?@        �       �                 pf�@ �#�Ѵ�?            �E@       ������������������������       �                     9@        �       �                 �|�=@�����H�?             2@       �       �                  sW@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 @3�@�_�s���?|            @i@        �       �                   �=@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    @<$c*(��?w            `h@       �       �                   �0@`����e�?o            �f@        �       �                    �?������?
             .@       �       �                 �̌!@d}h���?	             ,@        ������������������������       �                     @        �       �                    )@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �*@�+Ĺ+�?e            �d@       �       �                     @���2j��??            �Y@        �       �                    �?$G$n��?            �B@       �       �                 `fF)@؇���X�?            �A@        ������������������������       �        	             .@        �       �                    @@      �?             4@        ������������������������       �                     "@        �       �                   �F@�eP*L��?             &@        �       �                    C@r�q��?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �2@���Ls�?*            @P@        �       �                   �1@�z�G��?             $@        ������������������������       �                     @        �       �                 ��Y @      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�1�`jg�?&            �K@       �       �                 �|Y=@�X�<ݺ?%             K@        �       �                   �:@�t����?             1@       ������������������������       �        
             (@        �       �                 0S%"@���Q��?             @        ������������������������       �                     �?        �       �                 ���"@      �?             @        ������������������������       �                     �?        �       �                   �<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �"@�?�|�?            �B@       ������������������������       �                    �@@        �       �                 �|�=@      �?             @        ������������������������       �                      @        �       �                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�>@     ��?&             P@        �       �                 03�6@Pa�	�?            �@@       ������������������������       �                     :@        �       �                 03�7@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ?@        ������������������������       �                     ,@        �       �                    �?      �?              @       �       �                    ;@z�G�z�?             @        ������������������������       �                      @        �       �                    >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������v�S(��?��X��?�@ �?��~����?e�e��?�&�&�?��{a�?�{a���?F]t�E�?]t�E�?�a�a�?z��y���?�i�i�?\��[���?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?{�G�z�?���Q��?      �?                      �?      �?                      �?9��8���?�8��8��?�a�a�?�<��<��?�������?ZZZZZZ�?UUUUUU�?UUUUUU�?              �?]t�E�?F]t�E�?�������?UUUUUU�?              �?      �?              �?                      �?�{a���?a����?              �?�������?333333�?              �?      �?        �<ݚ�?���Hx�?��RJ)��?k���Zk�?UUUUUU�?UUUUUU�?              �?      �?        'u_[�?[4���?              �?|���?|���?�$I�$I�?�m۶m��?      �?      �?              �?      �?              �?      �?              �?      �?                      �?�5��P�?y�5���?      �?      �?�������?�������?      �?                      �?      �?        ]t�E�?t�E]t�?�$I�$I�?۶m۶m�?              �?      �?              �?              �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���͉�?�������?��Zk���?�RJ)���?UUUUUU�?�������?      �?      �?      �?                      �?              �?[�~�u��?J��/�?-n����?�#{���?�؉�؉�?�;�;�?UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?333333�?�������?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?F]t�E�?/�袋.�?              �?      �?      �?      �?                      �?�!5�x+�?�x+�R�?      �?      �?      �?                      �?/����?և���X�?      �?        ��L���?L�Ϻ��?------�?�������?�s�9��?�c�1Ƹ?�������?�?�q�q�?�q�q�?      �?        9��8���?�q�q�?      �?        �m۶m��?�$I�$I�?333333�?�������?      �?              �?                      �?      �?                      �?      �?        D8�C8��?�����?����!�?�琚`��?ڨ�l�w�?L� &W�?UUUUUU�?UUUUUU�?I�$I�$�?۶m۶m�?ffffff�?333333�?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?��Moz��?Y�B��?      �?              �?      �?      �?      �?      �?              �?      �?      �?      �?      �?              �?      �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?�������?333333�?      �?              �?      �?              �?      �?      �?      �?                      �?              �?,�����?�Σ�)�?gZ{���?e�,%l��?�]?[��?�F�tj�?
ףp=
�?���Q��?�Mozӛ�?d!Y�B�?      �?        �.�袋�?F]t�E�?      �?              �?      �?�������?�?�؉�؉�?;�;��?      �?              �?        ���8+�?�cj`?*�Y7�"�?к����?      �?        �/����?�}A_Ч?      �?        �q�q�?�q�q�?/�袋.�?F]t�E�?              �?      �?              �?              �?              �?        ��g����?Q`ҩy�?�$I�$I�?۶m۶m�?      �?                      �?��9��9�?�1�1�?jc��?X�s��C�?�?wwwwww�?۶m۶m�?I�$I�$�?              �?333333�?ffffff�?              �?      �?              �?        (፦ί�?���ˊ��?�������?�������?к����?���L�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?        t�E]t�?]t�E�?UUUUUU�?�������?              �?      �?      �?      �?              �?        �����?z�z��?ffffff�?333333�?      �?              �?      �?              �?      �?        A��)A�?�־a�?��8��8�?�q�q�?<<<<<<�?�?      �?        333333�?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?*�Y7�"�?к����?      �?              �?      �?      �?              �?      �?              �?      �?              �?             ��?      �?|���?|���?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?              �?              �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJt�mUhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM	hjh))��}�(h,h/h0M	��h2h3h4hph<�h=Kub������       ^                    �?<C�`��?�           8�@               %                     @�&��b�?�            �m@                                   �?d���i�?W            �a@                                  �?(�5�f��?-            �S@        ������������������������       �                    �A@                                   �?t��ճC�?             F@       ������������������������       �                     :@               	                    �?r�q��?
             2@       ������������������������       �                     *@        
                            @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @               $                    �?��� ��?*             O@                                 �B@�<ݚ�?             B@                                  �?HP�s��?             9@        ������������������������       �                     @                                  �;@ףp=
�?             4@                                  �6@�<ݚ�?             "@       ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                     �?                                  �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             &@               !                    �?�eP*L��?             &@                                  �*@�q�q�?             @                                  F@�q�q�?             @        ������������������������       �                     �?                                  �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        "       #                   �E@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        &       ]                   @B@D�]�+��?D            �X@       '       V                  ��8@(����7�?>            @V@       (       U                    @p9W��S�?5             S@       )       >                   �<@�M;q��?4            �R@       *       +                    @�&!��?            �E@        ������������������������       �                     @        ,       1                 ��,#@)O���?             B@        -       .                    �?r�q��?             2@        ������������������������       �                     @        /       0                   �7@�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @        2       9                    �?�<ݚ�?             2@        3       8                    �?���Q��?             @       4       5                 �&�)@�q�q�?             @        ������������������������       �                     �?        6       7                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        :       =                    �?8�Z$���?             *@        ;       <                   �8@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ?       T                    �?     ��?             @@       @       A                 �|Y=@д>��C�?             =@        ������������������������       �                      @        B       S                    �?�+$�jP�?             ;@       C       R                    �?H%u��?             9@       D       E                    �?��2(&�?             6@        ������������������������       �                     �?        F       M                   �>@�����?             5@       G       L                 �|�=@�IєX�?             1@       H       I                  ��@��S�ۿ?             .@        ������������������������       �                     @        J       K                 �̌'@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        N       Q                   �@@      �?             @       O       P                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        W       X                    �?$�q-�?	             *@        ������������������������       �                     �?        Y       Z                 ��T?@�8��8��?             (@        ������������������������       �                     @        [       \                 ��p@@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        _       �                    �?��lJ���?#           �}@       `       �                    �?��#�@��?�            �x@        a       p                     @4�{Y���?7            �T@        b       o                 p�w@�����H�?             ;@       c       d                    C@$�q-�?             :@       ������������������������       �        
             ,@        e       j                 p�i@@r�q��?             (@        f       i                     �?�q�q�?             @       g       h                  �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        k       l                    �?�����H�?             "@        ������������������������       �                     @        m       n                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        q       �                    �?����>4�?%             L@       r       u                   �5@�iʫ{�?#            �J@        s       t                 �y.@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        v       �                    �?      �?              H@       w       �                 ��$1@؇���X�?             E@       x       y                 ���@,���i�?            �D@        ������������������������       �                     "@        z                        �|Y=@     ��?             @@        {       |                    �?�q�q�?             @        ������������������������       �                      @        }       ~                  ��@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?ȵHPS!�?             :@        �       �                   @@����X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        �       �                 ���@�}�+r��?             3@        ������������������������       �                     @        �       �                   @'@��S�ۿ?             .@       �       �                 X�I@@4և���?             ,@       ������������������������       ��8��8��?             (@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                  �v6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?T>D5j�?�            �s@       �       �                 `fF:@���z�k�?�            Ps@       �       �                     @h�U���?�             o@        �       �                 `f�)@�k~X��?(             R@        ������������������������       �                     =@        �       �                   �*@ qP��B�?            �E@        �       �                   �C@�}�+r��?             3@       ������������������������       �                     0@        �       �                    G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        �       �                 �|�=@�O2�J�?r             f@       �       �                   �0@@A��q�?T            �`@        �       �                 �̌!@z�G�z�?             @       ������������������������       �      �?              @        ������������������������       �                     @        �       �                    �?0�ޤ��?Q            @`@       �       �                   �:@�(\����?L             ^@       ������������������������       �        -             S@        �       �                 0S%"@t��ճC�?             F@       �       �                 ��) @ףp=
�?             >@       �       �                 �?$@ 7���B�?             ;@        �       �                 ��,@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        �       �                 pf� @�q�q�?             @        ������������������������       �                     �?        �       �                 �|Y<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                     $@        �       �                   @@@؇���X�?             E@        �       �                    �?�q�q�?             (@       �       �                   �?@�eP*L��?             &@        �       �                   �>@�q�q�?             @       �       �                 �̌!@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �@���Q��?             @        ������������������������       �                     �?        �       �                 �?�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                 �?�@(;L]n�?             >@       ������������������������       �                     2@        �       �                   �D@�8��8��?             (@       �       �                   �B@      �?              @        ������������������������       �                     @        �       �                 ��	0@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     @d��0u��?$             N@       �       �                   �>@���dQ'�?!            �L@        �       �                    K@      �?             8@       �       �                   �<@@�0�!��?
             1@        ������������������������       �                     @        �       �                   @>@���!pc�?             &@       �       �                 �|�?@      �?              @        �       �                 �|Y=@      �?             @        ������������������������       �                     �?        �       �                 `fF<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 `fF<@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     �?6YE�t�?            �@@       �       �                 ��9L@     ��?             @@       �       �                    �?HP�s��?             9@       �       �                 ��yC@��S�ۿ?	             .@       �       �                 �|�<@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   @B@ףp=
�?             $@        ������������������������       �                     @        �       �                    G@r�q��?             @       �       �                  x#J@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 `f�N@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�r*e���?*            �R@        �       �                     @�8��8��?             (@       ������������������������       �                      @        �       �                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          �?r֛w���?#             O@       �                          �?�ՙ/�?             E@       �                        �y�/@^H���+�?            �B@        �       �                 ���"@�	j*D�?             *@        ������������������������       �                     @        �       �                 X�lA@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?                                 �?r�q��?             8@                                �B@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@                                 6@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     4@        �*       h�h))��}�(h,h/h0M	KK��h2h3h4hVh<�h=Kub�������������܍�W�?/�F�JP�?WAm���?��d~��?P$�Ҽ��?v{�e��?�&��jq�?�=Q���?              �?t�E]t�?�E]t��?              �?UUUUUU�?�������?              �?333333�?�������?      �?                      �?�B!��?�{����?�q�q�?9��8���?{�G�z�?q=
ףp�?              �?�������?�������?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�������?�������?              �?      �?                      �?/����?}h����?�9�as�?<��x��?l(�����?�k(����?ƒ_,���?�6�i��?S֔5eM�?֔5eMY�?              �?��8��8�?9��8���?UUUUUU�?�������?              �?�؉�؉�?ى�؉��?              �?      �?        9��8���?�q�q�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        ;�;��?;�;��?      �?      �?      �?                      �?      �?              �?      �?|a���?a���{�?              �?B{	�%��?/�����?���Q��?)\���(�?t�E]t�?��.���?      �?        �a�a�?=��<���?�?�?�?�������?              �?      �?      �?      �?                      �?              �?      �?      �?      �?      �?              �?      �?                      �?              �?      �?                      �?              �?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?              �?      �?              �?        �"h8���?'u_[�?�+2_�8�?�n-;�?�b��7��?4u~�!��?�q�q�?�q�q�?�؉�؉�?;�;��?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?n۶m۶�?I�$I�$�?
�[���?�琚`��?�������?333333�?              �?      �?              �?      �?۶m۶m�?�$I�$I�?�����?8��18�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?��N��N�?�؉�؉�?�m۶m��?�$I�$I�?      �?      �?      �?        �5��P�?(�����?      �?        �������?�?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?]ʥ\ʥ�?���Ѻ?���O ��?ch���V�?�����?��"NT��?�8��8��?�q�q�?      �?        ��}A�?�}A_З?�5��P�?(�����?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �v�,1�?k��2�?��)F�?t��:W�?�������?�������?      �?      �?      �?        /�B/�B�?z�z��?333333�?�������?      �?        �E]t��?t�E]t�?�������?�������?	�%����?h/�����?�������?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?              �?        ۶m۶m�?�$I�$I�?�������?�������?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?        DDDDDD�?wwwwww�?ZLg1���?Lg1��t�?      �?      �?�������?ZZZZZZ�?              �?t�E]t�?F]t�E�?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?۶m۶m�?�$I�$I�?      �?                      �?'�l��&�?e�M6�d�?      �?      �?q=
ףp�?{�G�z�?�������?�?۶m۶m�?�$I�$I�?              �?      �?              �?        �������?�������?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        0E>�S�?�u�)�Y�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        ���{��?�B!��?�<��<��?�a�a�?L�Ϻ��?�g�`�|�?;�;��?vb'vb'�?      �?        �������?�������?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?333333�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJc��hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM?hjh))��}�(h,h/h0M?��h2h3h4hph<�h=Kub������                        �Q��?ʡ�;S��?�           8�@        ������������������������       �                     "@               L                    �?����f��?�           ��@               +                     @�E�9��?]            `d@                                 �7@��}����?9            �X@                                  �6@�}�+r��?             3@       ������������������������       �                     *@               	                    �?r�q��?             @        ������������������������       �                     @        
                        �ܙC@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               (                     �?��Q��?.             T@              '                    �?.}Z*�?*            �Q@                                �>@�#��ؒ�?(            @Q@                                ��2>@�C��2(�?             &@                               ���<@z�G�z�?             @        ������������������������       �                      @                                X��@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �?�BbΊ�?!             M@       ������������������������       �                     ?@               "                 p"�X@X�<ݚ�?             ;@              !                    �?     ��?
             0@                               `f�A@X�<ݚ�?             "@        ������������������������       �                     @                                8�VQ@r�q��?             @       ������������������������       �                     @                                  �}S@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        #       &                    �?�C��2(�?             &@       $       %                 �̾w@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        )       *                    �?�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ,       I                 ��3@     ��?$             P@       -       <                 pF�#@^l��[B�?              M@       .       1                   �6@�S����?             C@        /       0                 ��y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        2       ;                 �|�=@      �?             @@       3       4                    �?      �?             0@        ������������������������       �                     �?        5       6                 ���@��S�ۿ?
             .@        ������������������������       �                     @        7       :                   @@ףp=
�?             $@       8       9                 �|=@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     0@        =       B                    �?��Q��?
             4@        >       ?                 0C1@�����H�?             "@        ������������������������       �                     @        @       A                   �2@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        C       D                    �?�eP*L��?             &@        ������������������������       �                     @        E       F                    7@؇���X�?             @        ������������������������       �                     @        G       H                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        J       K                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        M       �                     @8��X��?b           ؀@        N       e                    ,@�{���?�            `m@        O       \                    �?(���X�?)            @Q@        P       S                 ���&@z�G�z�?
             4@        Q       R                   �J@�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @        T       U                 ��Y)@؇���X�?             @        ������������������������       �                     �?        V       [                    D@r�q��?             @       W       Z                    �?�q�q�?             @       X       Y                    B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ]       d                    �?Hm_!'1�?            �H@       ^       _                    �?���}<S�?             G@        ������������������������       �                     �?        `       a                   �@@�:�^���?            �F@       ������������������������       �                     6@        b       c                   @A@�㙢�c�?             7@        ������������������������       ��q�q�?             @        ������������������������       �        	             1@        ������������������������       �                     @        f       �                    �?@K����?k            �d@       g       �                 `��R@l��[B��?I             ]@       h       �                   �G@� �	��?>             Y@       i       �                   �F@*-ڋ�p�?/            @S@       j       k                   �7@և���X�?)            �Q@        ������������������������       �                     @        l       �                     �?�G��l��?&            �O@       m       |                  x#J@�G��l��?             E@       n       o                    �?�n_Y�K�?             :@        ������������������������       �                     �?        p       u                 �|�<@��H�}�?             9@        q       r                   �;@      �?             @        ������������������������       �                     �?        s       t                 `f�D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        v       w                   @@@����X�?             5@       ������������������������       �                     "@        x       {                    �?      �?             (@       y       z                    D@�q�q�?             "@        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        }       ~                    �?      �?	             0@        ������������������������       �                     @               �                 `�iJ@���Q��?             $@        ������������������������       �                      @        �       �                    A@      �?              @       �       �                    7@�q�q�?             @        ������������������������       �                     �?        �       �                    <@z�G�z�?             @        ������������������������       �                      @        �       �                 `f�N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�ՙ/�?             5@        ������������������������       �                     @        �       �                   �E@��.k���?             1@       �       �                    �?��S���?
             .@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �J@�û��|�?             7@        �       �                 �D�J@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        �       �                    �?���|���?             &@        ������������������������       �                     @        �       �                 `fF<@      �?              @       ������������������������       �                     @        �       �                  )?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �C@      �?             0@       �       �                 �|�=@�����H�?             "@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?և���X�?             @        ������������������������       �                     @        �       �                   �G@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?j�q����?"             I@       �       �                    �?�(\����?             D@       ������������������������       �                     7@        �       �                    �?�IєX�?             1@        ������������������������       �                     @        �       �                 ��[@�C��2(�?             &@       ������������������������       �                     @        �       �                     @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        �       �                 �Cj]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    :@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       2                   @b_j�l�?�             s@       �       �                    @��0p'��?�            �p@        ������������������������       �                     @        �       �                    �?�Y����?�            �p@        �       �                 ��Y7@Υf���?)            �N@       �       �                    �?�û��|�?!             G@        �       �                    �?$�q-�?
             *@       �       �                 �|�9@ףp=
�?             $@        ������������������������       �                     �?        �       �                 ���@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    3@�'�=z��?            �@@        ������������������������       �                     @        �       �                   �.@*;L]n�?             >@       �       �                 ���@���!pc�?             6@        ������������������������       �                      @        �       �                   �9@z�G�z�?             4@        ������������������������       �                     $@        �       �                    ;@���Q��?             $@        ������������������������       �                      @        �       �                 ��n @      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                  SE"@�q�q�?             @        ������������������������       �                     �?        �       �                   &@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                 03�1@؇���X�?             @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�r����?             .@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @$�q-�?             *@        ������������������������       �                     @        �       �                   �C@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���}<S�?�            �i@        �       �                 �|Y=@�㙢�c�?             7@        �       �                  ��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?ףp=
�?             4@       �       �                    �?�KM�]�?             3@       �       �                    �?�X�<ݺ?             2@       �       �                  s�@@4և���?             ,@        ������������������������       �                     @        �       �                 X��A@�C��2(�?	             &@       �       �                   @'@�����H�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �                         �7@�c:��?x             g@        �                         �2@ _�@�Y�?%             M@        �       �                   �1@�}�+r��?             3@       ������������������������       �                     &@        �                          �?      �?              @       �                          �?r�q��?             @                              ���@z�G�z�?             @        ������������������������       �                     @                              ��Y @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �C@              +                  @@@|�(��?S            �_@       	      "                �|�=@PN��T'�?7            @T@       
                      ��) @�θV�?/            @Q@                                �?�nkK�?              G@                               @8@ �#�Ѵ�?            �E@                                �@���Q��?             @                              �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     C@        ������������������������       �                     @              !                   �?��<b���?             7@                                (@     ��?             0@                                �<@      �?              @                                �;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                              �|Y=@      �?             @        ������������������������       �                      @                              pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        #      &                �̌!@�q�q�?             (@       $      %                  �@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        '      (                ��Y)@z�G�z�?             @        ������������������������       �                     @        )      *                �!B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ,      1                  �C@����?�?            �F@       -      0                @3�@���7�?             6@        .      /                  @C@؇���X�?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �        	             .@        ������������������������       �                     7@        3      4                   �?�FVQ&�?            �@@        ������������������������       �        
             0@        5      8                   �?�t����?             1@       6      7                ���1@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        9      >                pf�C@      �?              @        :      ;                   @      �?             @        ������������������������       �                     �?        <      =                   @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M?KK��h2h3h4hVh<�h=Kub������������N���I5�?d�~`l��?              �?zG"Ϝw�?q�a��?�E:i�?�r��bK�?P�W
���?X
����?(�����?�5��P�?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?ffffff�?�������?�
��V�?�z2~���?s��\;0�?F��Q�g�?]t�E�?F]t�E�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ���=��?�{a��?              �?r�q��?�q�q�?      �?      �?r�q��?�q�q�?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?]t�E�?F]t�E�?�������?UUUUUU�?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?�=�����?��=���?(������?^Cy�5�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?              �?�������?�?      �?        �������?�������?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?        �������?ffffff�?�q�q�?�q�q�?      �?              �?      �?      �?                      �?]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?UUUUUU�?�������?      �?                      �?L3��@��?i��~/�?sB�n�?{��#��?l�ځ��?)�3J���?�������?�������?�؉�؉�?ى�؉��?              �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?Y�Cc�?9/���?ӛ���7�?d!Y�B�?      �?        }�'}�'�?l�l��?      �?        �7��Mo�?d!Y�B�?UUUUUU�?UUUUUU�?      �?              �?        �b��7��?�ί=��?���=��?GX�i���?�Q����?)\���(�??!��O��?��cj`��?�$I�$I�?۶m۶m�?      �?        1�0��?��y��y�?��y��y�?1�0��?;�;��?ى�؉��?              �?{�G�z�?
ףp=
�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?              �?�������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �<��<��?�a�a�?      �?        �������?�?�������?�?              �?      �?              �?              �?        ��,d!�?8��Moz�?UUUUUU�?�������?              �?      �?        ]t�E]�?F]t�E�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?
ףp=
�?=
ףp=�?�������?333333�?              �?�?�?              �?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?�������?�������?      �?      �?              �?      �?              �?      �?              �?      �?        ����k�?�5��P�?�&�U��?e��?              �?��¯�D�?���@���?i�>�%C�?.�u�y�?��,d!�?8��Moz�?;�;��?�؉�؉�?�������?�������?              �?�q�q�?�q�q�?      �?                      �?              �?|��|�?|���?              �?""""""�?�������?F]t�E�?t�E]t�?              �?�������?�������?      �?        333333�?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?      �?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?�������?�?      �?      �?      �?                      �?�؉�؉�?;�;��?      �?        ۶m۶m�?�$I�$I�?              �?      �?        ӛ���7�?d!Y�B�?�7��Mo�?d!Y�B�?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?�k(���?(�����?��8��8�?�q�q�?n۶m۶�?�$I�$I�?      �?        ]t�E�?F]t�E�?�q�q�?�q�q�?      �?      �?      �?              �?              �?                      �?      �?        Y�B���?8��Moz�?#,�4�r�?�{a���?�5��P�?(�����?      �?              �?      �?�������?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?              �?              �?              �?        -˲,˲�?��i��i�?&���^B�?h/�����?̵s���?�Q�g���?�Mozӛ�?d!Y�B�?�/����?�}A_Ч?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        ��,d!�?��Moz��?      �?      �?      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?              �?      �?              �?        �������?�������?۶m۶m�?�$I�$I�?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?��I��I�?l�l��?�.�袋�?F]t�E�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?              �?        >����?|���?      �?        <<<<<<�?�?�q�q�?�q�q�?              �?      �?              �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg�$hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM?hjh))��}�(h,h/h0M?��h2h3h4hph<�h=Kub������       h                    �?|��;;��?�           8�@               g                    @C��3�?�            @o@              6                   �;@�Ee@���?�            �n@                                    @J��D��?D             [@                                    �? i���t�?            �H@                                   �?P���Q�?             4@       ������������������������       �                     *@               	                    �?؇���X�?             @       ������������������������       �                     @        
                           )@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �7@\-��p�?             =@       ������������������������       �                     4@                                   �?X�<ݚ�?             "@        ������������������������       �                     �?                                   �?      �?              @                                  �9@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                  �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               -                   �3@�m����?%            �M@                               ��*@�t����?             A@        ������������������������       �                     2@               (                    @      �?             0@              '                 ��*4@���!pc�?
             &@              $                    �?և���X�?             @                                  �?      �?             @        ������������������������       �                     �?                #                    �?�q�q�?             @       !       "                    (@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        %       &                  �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        )       ,                    @���Q��?             @       *       +                 ��T?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        .       /                 pf&@�+e�X�?             9@        ������������������������       �                     @        0       5                 pf� @P���Q�?	             4@        1       4                    �?�����H�?             "@       2       3                   �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        7       D                 `f�$@0Lj����?Y             a@        8       C                    �?���Q��?             4@       9       B                    A@      �?             0@       :       ?                    �?؇���X�?             ,@       ;       >                 ���@�C��2(�?	             &@        <       =                 �Y�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        @       A                 ��; @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        E       P                     @�q3�M��?J             ]@       F       G                     �?��f�{��?7            �U@       ������������������������       �                     G@        H       I                    9@�(\����?             D@       ������������������������       �                     :@        J       O                    �?@4և���?
             ,@       K       L                    �?      �?              @        ������������������������       �                      @        M       N                    D@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        Q       Z                    �?�q�q�?             >@       R       S                    �?�}�+r��?
             3@        ������������������������       �                     "@        T       Y                     @ףp=
�?             $@       U       X                 ���.@      �?              @        V       W                 ���*@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        [       b                   �>@"pc�
�?	             &@       \       a                 `v�6@      �?              @        ]       ^                 �|�<@      �?             @        ������������������������       �                     �?        _       `                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        c       d                 hV}1@�q�q�?             @        ������������������������       �                     �?        e       f                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        i       �                     �?`�N�?           �|@        j       �                    �?��_����?=            �[@       k       �                 �̾w@$��m��?:             Z@       l       �                    �?�g��@(�?9            @Y@       m       �                   �H@�q�q�?3            �V@       n       o                   �9@4���C�?&            �P@        ������������������������       �                     @        p       �                  �>@N1���?$            �N@        q       r                   �;@��Q��?             4@        ������������������������       �                      @        s       |                 ���<@b�2�tk�?             2@       t       u                    @@      �?             (@        ������������������������       �                     @        v       w                 03k:@      �?              @        ������������������������       �                     �?        x       y                   �C@����X�?             @        ������������������������       �                     @        z       {                   @G@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        }       �                   @>@r�q��?             @       ~                        �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 �!�I@��]�T��?            �D@        �       �                 �|�<@�����H�?
             2@        �       �                 `f�D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��S�ۿ?             .@        �       �                  �>@z�G�z�?             @        ������������������������       �                      @        �       �                    C@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �8@\X��t�?             7@        ������������������������       �                     @        �       �                    �?�����?
             3@        ������������������������       �                     @        �       �                 �w|c@և���X�?             ,@       �       �                   �D@���!pc�?             &@       �       �                 03�S@z�G�z�?             $@       �       �                 `f�N@����X�?             @       �       �                 `f�K@r�q��?             @       �       �                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���=@�8��8��?             8@        ������������������������       �                     (@        �       �                   �R@r�q��?             (@       �       �                    �?�C��2(�?             &@        ������������������������       �                     @        �       �                   �I@r�q��?             @        ������������������������       �                     @        �       �                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���!pc�?             &@       �       �                   �7@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    /@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�:pΈ��?�            �u@        �       �                     @      �?!             H@        ������������������������       �                     $@        �       �                    �?�����?             C@       �       �                 �|Y=@V�a�� �?             =@        �       �                    �?�eP*L��?             &@       �       �                 ��y@���Q��?             $@        ������������������������       �                      @        �       �                    /@      �?              @        ������������������������       �                      @        �       �                   �6@�q�q�?             @        ������������������������       �                     @        �       �                   �<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y?@�X�<ݺ?             2@       �       �                   @@�C��2(�?	             &@       �       �                 ���@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �x"@�q�q�?             "@        ������������������������       �                     �?        �       �                 �&�)@      �?              @        ������������������������       �                     @        �       �                    7@      �?             @        ������������������������       �                     �?        �       �                 �|Y<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       .                   �?�4�����?�            �r@       �       '                0��D@��F!�?�            �l@       �       �                    )@<\����?�            �k@        ������������������������       �                     @        �       �                     @��n5V�?�            `k@        �       �                    5@(;L]n�?%             N@        �       �                    &@      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                   @@@ pƵHP�?!             J@        ������������������������       �                     9@        �       �                   �*@ 7���B�?             ;@       �       �                   @A@�IєX�?             1@        ������������������������       ��q�q�?             @        ������������������������       �        	             ,@        ������������������������       �                     $@        �       �                    �?�J��_��?h            �c@        �       �                 �|Y;@@4և���?	             ,@        ������������������������       �                     �?        �       �                 X��A@$�q-�?             *@       �       �                 ���@�8��8��?             (@        ������������������������       �                     @        �       �                 ��(@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �0@������?_             b@        �       �                 pFD!@�q�q�?             @        �       �                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       &                   �?��*��?[            `a@       �                       �|Y>@�<_���?Z             a@       �                       @3�@(a��䛼?E            @Y@       �       �                    7@h�����?%             L@        ������������������������       �                     2@        �                       �?$@�}�+r��?             C@        �       �                   �8@�����H�?             2@        �       �                 �&b@r�q��?             @        ������������������������       �                     @        �       �                 `fF@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                        ���@�8��8��?	             (@       ������������������������       �                     "@                              �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     4@              
                  �:@�:�^���?             �F@              	                0S5 @���7�?             6@                                �3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@                                �;@�LQ�1	�?             7@        ������������������������       �                     �?                              ��) @�C��2(�?             6@        ������������������������       �                     $@                                �<@r�q��?	             (@        ������������������������       �                     @                              pf� @      �?              @        ������������������������       �                     �?                              ��)"@؇���X�?             @        ������������������������       �                     @                              �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @              !                  @@@4?,R��?             B@                                �?@�q�q�?             "@                              pff@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?                              P�@      �?             @        ������������������������       �                     �?                               ��I @�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        "      #                �?�@�>����?             ;@       ������������������������       �        
             2@        $      %                @3�@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        (      )                  �7@և���X�?             @        ������������������������       �                      @        *      +                   ;@z�G�z�?             @        ������������������������       �                     @        ,      -                   >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        /      :                   �?��W��?-            @R@       0      5                    @r�qG�?             H@        1      2                  �3@8�A�0��?             6@        ������������������������       �                     @        3      4                   0@������?             1@        ������������������������       �                     @        ������������������������       �        	             *@        6      7                   �?8�Z$���?             :@        ������������������������       �                     @        8      9                   )@�㙢�c�?             7@        ������������������������       �                     @        ������������������������       �                     3@        ;      >                    @`2U0*��?             9@        <      =                  @9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        �*       h�h))��}�(h,h/h0M?KK��h2h3h4hVh<�h=Kub������������|d�_Z�?�7s@K�?h��|?5�?��� �r�?q�����?�����?_B{	�%�?�^B{	��?����X�?/�����?�������?ffffff�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?�{a���?a����?              �?�q�q�?r�q��?              �?      �?      �?�������?333333�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �V'u�?��}ylE�?�������?�������?              �?      �?      �?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?333333�?      �?      �?      �?                      �?      �?        R���Q�?���Q��?              �?ffffff�?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?�������?333333�?      �?      �?�$I�$I�?۶m۶m�?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �i��F�?�rO#,��?�}A_Ї?������?              �?�������?333333�?              �?�$I�$I�?n۶m۶�?      �?      �?              �?UUUUUU�?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?(�����?�5��P�?              �?�������?�������?      �?      �?      �?      �?              �?      �?                      �?              �?/�袋.�?F]t�E�?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        !�]����?}��29��?�B�I .�?<zel���?�N��N��?vb'vb'�?���g��?���(0��?UUUUUU�?UUUUUU�?m��&�l�?'�l��&�?      �?        �:ڼO�?�}�K�`�?ffffff�?�������?              �?9��8���?�8��8��?      �?      �?      �?              �?      �?              �?�$I�$I�?�m۶m��?              �?      �?      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?KԮD�J�?jW�v%j�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?        �������?�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ��Moz��?!Y�B�?      �?        ^Cy�5�?Q^Cy��?              �?۶m۶m�?�$I�$I�?t�E]t�?F]t�E�?�������?�������?�$I�$I�?�m۶m��?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?]t�E�?F]t�E�?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?                      �?F]t�E�?t�E]t�?ffffff�?333333�?              �?      �?              �?                      �?�$I�$I�?�m۶m��?              �?      �?        ��Q���?�Q����?      �?      �?      �?        Q^Cy��?^Cy�5�?��{a�?a���{�?t�E]t�?]t�E�?333333�?�������?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?��8��8�?�q�q�?]t�E�?F]t�E�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?aQ�(X�?�t}�>]�?یZ9��?'�+�7��?.Ԝ�B�?�^���?              �?��_j��?@+���?�������?�?      �?      �?      �?      �?      �?        'vb'vb�?;�;��?      �?        	�%����?h/�����?�?�?UUUUUU�?UUUUUU�?      �?              �?        d�^�.�?�%w��?n۶m۶�?�$I�$I�?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?      �?      �?              �?        ��y�!�?C:o1��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        4,�T�w�?c�>ZMB�?p�h�?n�?ܺ���?��~�X�?�F�tj�?�m۶m��?�$I�$I�?      �?        �5��P�?(�����?�q�q�?�q�q�?�������?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?        }�'}�'�?l�l��?�.�袋�?F]t�E�?�������?�������?              �?      �?              �?        ��Moz��?Y�B��?              �?]t�E�?F]t�E�?      �?        �������?UUUUUU�?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        �8��8��?r�q��?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        �Kh/��?h/�����?      �?        9��8���?�q�q�?              �?      �?              �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?      �?      �?                      �?ϝ;w���?Ĉ#F��?UUUUUU�?UUUUUU�?颋.���?/�袋.�?              �?xxxxxx�?�?              �?      �?        ;�;��?;�;��?      �?        �7��Mo�?d!Y�B�?              �?      �?        ���Q��?{�G�z�?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�>D5hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������                           @��ҴҰ�?�           8�@                                   @b�h�d.�?            �A@                               �-]@h�����?             <@       ������������������������       �                     :@                                �(\�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                ���A@����X�?             @       	       
                 ��T?@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               f                    �?*$9	��?�            �@               W                    �?>���Rp�?�             m@                                   @�������?�            `j@                               03�=@0x�!���?L            �]@                                   �?l�b�G��?$            �L@                               ���;@���}<S�?             G@                                  �? qP��B�?            �E@        ������������������������       �                     @                                  �;@�?�|�?            �B@                                  �9@�8��8��?             (@       ������������������������       �                     $@                                  �/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     9@        ������������������������       �                     @        ������������������������       �        	             &@        ������������������������       �        (             O@               V                   @C@<SvLB�?9             W@               !                    &@t�����?3             U@        ������������������������       �                     @        "       ?                    �?��Q���?2             T@       #       $                   �0@ �o_��?             I@        ������������������������       �                     @        %       >                    @p�v>��?            �G@       &       -                    �?8����?             G@        '       (                    �?��2(&�?             6@       ������������������������       �        
             1@        )       *                 ���&@���Q��?             @        ������������������������       �                      @        +       ,                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        .       9                 @33"@r�q��?             8@       /       8                 @3�@      �?
             0@       0       5                 �&B@��
ц��?             *@       1       4                   �7@r�q��?             @        2       3                    4@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        6       7                    ;@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        :       =                 ��&@      �?              @       ;       <                 �[$@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        @       A                 pF�%@*;L]n�?             >@        ������������������������       �                     @        B       U                   �@@�q�q�?             8@       C       T                    �?b�2�tk�?             2@       D       E                 �&�)@ҳ�wY;�?             1@        ������������������������       �                     @        F       K                    �?և���X�?             ,@        G       H                 �|6@      �?             @        ������������������������       �                      @        I       J                 P�h2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        L       Q                    �?�z�G��?             $@       M       N                    �?      �?              @        ������������������������       �                     @        O       P                 03�0@      �?             @        ������������������������       �                      @        ������������������������       �                      @        R       S                   �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        X       e                 �̾d@�ՙ/�?             5@       Y       ^                    �?������?             1@        Z       ]                    @      �?             @       [       \                 �|�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        _       `                   �6@$�q-�?             *@        ������������������������       �                      @        a       d                    �?z�G�z�?             @       b       c                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        g       �                  x#J@t�!ǐ��?           �{@       h       �                    �?ДX��?�            �y@        i       j                 ���@t�7��?$             O@        ������������������������       �                     (@        k       x                 �|Y=@H.�!���?             I@        l       s                 ��*@�q�q�?             .@        m       r                   @@X�<ݚ�?             "@       n       q                   @8@����X�?             @       o       p                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        t       u                 0C�<@r�q��?             @        ������������������������       �                     @        v       w                   �9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        y       �                    �?b�h�d.�?            �A@       z       �                    �?�r����?             >@       {       |                    A@؇���X�?             <@       ������������������������       �                     0@        }       ~                 `f�3@�q�q�?             (@        ������������������������       �                     @               �                    H@      �?              @       �       �                   �A@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     @���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                     �?H������?�            �u@        �       �                   �B@8�Z$���?             J@       �       �                 �|�<@r٣����?            �@@        ������������������������       �                     �?        �       �                   �J@     ��?             @@       �       �                   �G@R�}e�.�?             :@       �       �                   �B@�㙢�c�?             7@       �       �                    A@������?
             1@       �       �                 `fF<@     ��?	             0@       ������������������������       �                     &@        �       �                   �>@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             3@        �       �                   @A@��v�u�?�            `r@       �       �                    �?=�J�C�?�            �m@       �       �                     @`�a�?�            `i@        �       �                    @     ��?             @@        ������������������������       �                     @        �       �                    &@�+e�X�?             9@        ������������������������       ��q�q�?             @        �       �                 �|Y;@"pc�
�?             6@       ������������������������       �                     ,@        �       �                 �|�=@      �?              @        ������������������������       �                     @        �       �                    @@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        �       �                 �|�=@�� ND��?n            `e@       �       �                 ���@�O��e�?`            �b@        ������������������������       �                     ;@        �       �                   �3@4Qi0���?N            �^@        �       �                 0S5 @������?             1@        �       �                   �1@X�<ݚ�?             "@        ������������������������       �      �?             @        �       �                 �?�@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        �       �                   �:@�8�l��?C            �Z@        ������������������������       �                    �@@        �       �                 �?$@����1�?,            @R@        �       �                 ��@���N8�?             5@       �       �                 �|Y=@r�q��?	             2@        ������������������������       �                      @        ������������������������       �      �?             0@        ������������������������       ��q�q�?             @        �       �                 ��) @ ��WV�?!             J@       ������������������������       �                     C@        �       �                 ��)"@؇���X�?	             ,@        ������������������������       �                      @        ������������������������       �                     (@        �       �                   @@@���N8�?             5@       �       �                 ���!@�eP*L��?
             &@       �       �                   �>@�q�q�?	             "@        ������������������������       �                      @        �       �                   �?@և���X�?             @        �       �                 pff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �@���Q��?             @        ������������������������       �                     �?        �       �                 �?�@      �?             @        ������������������������       �                     �?        �       �                 ��I @�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?������?             B@       �       �                     @ ��WV�?             :@        ������������������������       �                     @        �       �                    7@���N8�?             5@        �       �                    �?�����H�?             "@        �       �                  s�@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �        	             $@        ������������������������       �        $            �K@        �       �                    �?*O���?             B@       �       �                   �E@�G��l��?             5@       �       �                 ���X@      �?             0@       �       �                     �?����X�?	             ,@       �       �                   �9@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                     @�q�q�?             @        ������������������������       �                     �?        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 @�:x@z�G�z�?	             .@       �       �                    �?$�q-�?             *@        �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �                  "&d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub���������������(�TL�?���Vg�?_�_��?;��:���?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?        �m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        �Z$���?:J�����?GX�i���?�i��F�?�Y����?�iP�z�?�5�5�?��~���?p�}��?�Gp��?d!Y�B�?ӛ���7�?�}A_З?��}A�?              �?к����?*�Y7�"�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?                      �?              �?���,d!�?�7��Mo�?�y��y��?�0�0�?      �?        �������?333333�?�Q����?
ףp=
�?              �?L� &W�?ڨ�l�w�?8��Moz�?d!Y�B�?t�E]t�?��.���?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?�;�;�?�؉�؉�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?�m۶m��?              �?      �?              �?              �?      �?      �?      �?              �?      �?                      �?              �?�������?""""""�?      �?        �������?�������?9��8���?�8��8��?�������?�������?              �?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?      �?                      �?333333�?ffffff�?      �?      �?              �?      �?      �?              �?      �?              �?      �?      �?                      �?      �?                      �?      �?        �<��<��?�a�a�?xxxxxx�?�?      �?      �?      �?      �?      �?                      �?              �?�؉�؉�?;�;��?      �?        �������?�������?      �?      �?              �?      �?              �?                      �?�@\�9	�?c��2��?�������?ZZZZZZ�?SJ)��R�?��Zk���?      �?        �(\����?)\���(�?UUUUUU�?UUUUUU�?r�q��?�q�q�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?;��:���?_�_��?�������?�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?�������?�������?              �?      �?              �?              �?        333333�?�������?      �?                      �?T���"�?]����?;�;��?;�;��?>���>�?|���?              �?      �?      �?'vb'vb�?�;�;�?�7��Mo�?d!Y�B�?xxxxxx�?�?      �?      �?      �?        �������?333333�?              �?      �?                      �?      �?                      �?      �?              �?        `��!�?e�J��?WAm���?J���Ϣ�?�^q2��?Ztl��?      �?      �?      �?        R���Q�?���Q��?UUUUUU�?UUUUUU�?/�袋.�?F]t�E�?      �?              �?      �?              �?�������?�������?      �?              �?      �?�_@�?@���?�t�@��?ƒ_,�Ų?      �?        #6�a#�?�On��?xxxxxx�?�?r�q��?�q�q�?      �?      �?333333�?�������?      �?              �?      �?      �?        �>����?�	�[��?      �?        �Ν;w��?Ĉ#F��?�a�a�?��y��y�?�������?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?O��N���?;�;��?      �?        ۶m۶m�?�$I�$I�?              �?      �?        �a�a�?��y��y�?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?333333�?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �q�q�?�q�q�?O��N���?;�;��?      �?        ��y��y�?�a�a�?�q�q�?�q�q�?      �?      �?      �?                      �?      �?              �?              �?              �?        �q�q�?�q�q�?1�0��?��y��y�?      �?      �?�$I�$I�?�m۶m��?F]t�E�?/�袋.�?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?        �������?�������?�؉�؉�?;�;��?�������?�������?      �?              �?      �?              �?      �?              �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���&hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       \                    �?"��p�?�           8�@                                    @6�I#r�?�             o@                                  �?���Z�?Y             a@        ������������������������       �                    �D@                                    �?p�qG�??             X@                                   �?P���Q�?             D@       ������������������������       �                     8@                                   �?      �?             0@       	       
                 ��1^@8�Z$���?             *@       ������������������������       �                     "@                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                  �J@�h����?$             L@                                  6@@3����?#             K@                                   �?�IєX�?             1@       ������������������������       �                     0@        ������������������������       �                     �?        ������������������������       �                    �B@        ������������������������       �                      @               K                 ���4@և���X�?H             \@              ,                 �̌@PN���?9            @V@               +                 X��B@�MI8d�?            �B@              *                    �?4?,R��?             B@              !                    �?��hJ,�?             A@                               �|Y8@�}�+r��?             3@        ������������������������       �                     @                                   �?@4և���?
             ,@        ������������������������       �                     �?                                 ���@$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        "       #                  s@������?             .@        ������������������������       �                     @        $       %                    4@�q�q�?             (@        ������������������������       �                     @        &       )                 pf�@�����H�?             "@        '       (                 �|Y:@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        -       6                 `f�%@
j*D>�?#             J@        .       /                    �?�S����?             3@        ������������������������       �                     �?        0       5                 @3�@�����H�?             2@        1       2                 �?�@����X�?             @        ������������������������       �                      @        3       4                   �9@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        7       @                    �?"pc�
�?            �@@        8       9                 P��+@�q�q�?             "@        ������������������������       �                     @        :       ;                 �?�-@      �?             @        ������������������������       �                      @        <       ?                    �?      �?             @       =       >                    3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        A       B                   �*@      �?             8@        ������������������������       �                     @        C       D                    .@@�0�!��?             1@        ������������������������       �                      @        E       F                    �?��S�ۿ?	             .@        ������������������������       �                     @        G       H                   @1@�C��2(�?             &@       ������������������������       �                     @        I       J                   �8@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        L       M                    �?�LQ�1	�?             7@        ������������������������       �                     �?        N       S                    @�C��2(�?             6@        O       P                    @�q�q�?             @        ������������������������       �                     �?        Q       R                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        T       U                 ��T?@�}�+r��?             3@       ������������������������       �                     $@        V       W                    �?�����H�?             "@        ������������������������       �                     @        X       [                    @r�q��?             @        Y       Z                 ��p@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ]       �                 03c4@F��ʁ�?           �|@       ^       q                    �?�KM�]�?�             s@        _       `                 =
�@�p ��?            �D@        ������������������������       �                     �?        a       b                    5@      �?             D@        ������������������������       �                      @        c       n                    �?     ��?             @@       d       m                 �� @8�Z$���?             :@       e       l                   @@���y4F�?             3@       f       i                 ���@�t����?             1@       g       h                 �|�9@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        j       k                 �|=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     @        o       p                 �|Y<@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        r       s                     �?X�g�Y��?�            pp@        ������������������������       �                     @        t       �                 �?�@�|K��2�?�             p@        u       �                    �?@\�*��?H            @]@       v       w                     @`����x�?F            �\@        ������������������������       �                     @        x       {                    �?���7�?C            �[@        y       z                 �|Y=@@4և���?             <@        ������������������������       �                      @        ������������������������       �                     :@        |       �                   �@Ћ����?5            �T@       }       �                 P�N@�1�`jg�?#            �K@       ~                           7@@9G��?            �H@        ������������������������       �        	             3@        �       �                 �&b@��S�ۿ?             >@        ������������������������       �                     $@        �       �                 ���@ףp=
�?             4@        ������������������������       �                     �?        �       �                 �|Y>@�}�+r��?             3@       �       �                 pf�@@4և���?	             ,@        ������������������������       �                      @        �       �                 �|�<@r�q��?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                    >@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ;@        ������������������������       �                     @        �       �                    �?��0{9�?\            �a@       �       �                   �2@(��R%��?U            �`@        �       �                   �0@X�Cc�?             ,@        �       �                 pFD!@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                 pf� @����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �:@POͳF��?N            �]@        �       �                 ���$@P�Lt�<�?             C@       ������������������������       �                     6@        �       �                    4@      �?             0@        �       �                   �'@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?PN��T'�?5            @T@       �       �                   @A@r�q��?0             R@       �       �                 @3�@      �?             F@        ������������������������       �                     @        �       �                 `fF)@z�G�z�?             D@       �       �                     @ףp=
�?             >@        ������������������������       �                     @        �       �                   �;@      �?             8@        ������������������������       �                     �?        �       �                 �|Y=@���}<S�?             7@        �       �                   �<@z�G�z�?             @        ������������������������       �                      @        �       �                 ���"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �y'"@�X�<ݺ?             2@       ������������������������       �        
             *@        �       �                 �|�=@z�G�z�?             @        ������������������������       �                      @        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     @���Q��?             $@       �       �                 �|�<@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�=@z�G�z�?             @        ������������������������       �                      @        �       �                    @@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 @3�@h�����?             <@        ������������������������       ��q�q�?             @        ������������������������       �                     9@        ������������������������       �                     "@        �       �                    �?      �?              @       �       �                    &@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �                            �?0h���b�?_            �c@       �       �                   �J@�E���?<            @X@       �       �                    �?yÏP�?2            �T@        �       �                   �8@     ��?             @@        ������������������������       �                     @        �       �                 p�w@��>4և�?             <@       �       �                    �?      �?             6@       �       �                 �|�;@ҳ�wY;�?
             1@        ������������������������       �                     @        �       �                   @@@��
ц��?             *@        �       �                 �|�=@r�q��?             @       �       �                 03SA@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �A@؇���X�?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �G@��H�}�?              I@       �       �                    �?���!pc�?             F@       �       �                   �>@�%^�?            �E@        �       �                    D@�z�G��?             $@       �       �                 �|�?@؇���X�?             @       �       �                 �|�<@      �?             @        ������������������������       �                      @        �       �                 `f�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                   �;@<���D�?            �@@        ������������������������       �                     �?        �       �                    �?     ��?             @@       �       �                 `f�D@ �q�q�?             8@        �       �                 �|�<@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        �       �                 03�S@      �?              @       �       �                    A@؇���X�?             @        �       �                    >@�q�q�?             @        ������������������������       �                     �?        �       �                   @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �R@��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?                                 �?��f/w�?#            �N@        ������������������������       �                     @                              ���4@�MWl��?!            �L@        ������������������������       �                     @                                 @�+$�jP�?             K@                                  @և���X�?             ,@        ������������������������       �                     @        ������������������������       �                      @        	                         �?ףp=
�?             D@        
                      0��D@������?             1@                                �?ףp=
�?             $@                              03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                              �|�>@և���X�?             @                             ��?P@z�G�z�?             @                                ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������J54v��?l�����?a2�>�?h3�?R0�?T{N���?�J���?              �?�������?UUUUUU�?�������?ffffff�?              �?      �?      �?;�;��?;�;��?              �?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?h/�����?���Kh�?�?�?              �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?B�P�"�?_��׽��?L�Ϻ��?��L���?r�q��?�8��8��?�������?KKKKKK�?(�����?�5��P�?              �?�$I�$I�?n۶m۶�?              �?;�;��?�؉�؉�?      �?                      �?�?wwwwww�?              �?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?      �?      �?              �?      �?                      �?              �?      �?        ;�;��?b'vb'v�?(������?^Cy�5�?              �?�q�q�?�q�q�?�m۶m��?�$I�$I�?      �?        333333�?�������?      �?                      �?      �?        F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?      �?      �?                      �?              �?      �?      �?              �?�������?ZZZZZZ�?      �?        �?�������?              �?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?��Moz��?Y�B��?              �?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�5��P�?(�����?      �?        �q�q�?�q�q�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        �����c�?(�Y�	q�?�k(���?(�����?Q��+Q�?��+Q��?              �?      �?      �?      �?              �?      �?;�;��?;�;��?6��P^C�?(������?<<<<<<�?�?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?              �?      �?              �?      �?        �������?UUUUUU�?      �?                      �?�p�$��?�x\�N�?      �?        2g�s��?sƜ1g̹?���?^�^�?��,����?Lg1��t�?      �?        �.�袋�?F]t�E�?n۶m۶�?�$I�$I�?              �?      �?        ԮD�J��?��+Q��?A��)A�?�־a�?������?9/���?      �?        �������?�?      �?        �������?�������?              �?�5��P�?(�����?n۶m۶�?�$I�$I�?      �?        �������?UUUUUU�?      �?              �?      �?      �?        �������?UUUUUU�?      �?                      �?      �?              �?        m�w6�;�?L� &W�?����N��?,�T�R�?%I�$I��?�m۶m��?�$I�$I�?۶m۶m�?      �?      �?      �?        �m۶m��?�$I�$I�?              �?      �?        ]�\��?e�e��?���k(�?(�����?      �?              �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?        &���^B�?h/�����?�������?UUUUUU�?      �?      �?              �?ffffff�?ffffff�?�������?�������?      �?              �?      �?              �?ӛ���7�?d!Y�B�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?��8��8�?�q�q�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?              �?      �?      �?      �?              �?      �?              �?        '��jq�?�g *��?tT����?W?���?W�v%jW�?Q��+Q�?      �?      �?      �?        I�$I�$�?۶m۶m�?      �?      �?�������?�������?              �?�؉�؉�?�;�;�?�������?UUUUUU�?      �?      �?              �?      �?              �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?                      �?{�G�z�?
ףp=
�?F]t�E�?t�E]t�?�}A_��?�}A_�?333333�?ffffff�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?|���?|���?              �?      �?      �?�������?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?              �?              �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?              �?              �?�������?�?      �?                      �?XG��).�?��!XG�?      �?        :��,���?�YLg1�?              �?/�����?B{	�%��?�$I�$I�?۶m۶m�?              �?      �?        �������?�������?xxxxxx�?�?�������?�������?      �?      �?              �?      �?              �?        �$I�$I�?۶m۶m�?�������?�������?      �?      �?              �?      �?              �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�EhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM?hjh))��}�(h,h/h0M?��h2h3h4hph<�h=Kub������       �                    �?>AU`�z�?�           8�@              /                    �?��\�#�?(           �}@                                ��4=@R�����?5             T@                                  �?���N8�?             E@                                X��B@      �?              @       ������������������������       �                     @        ������������������������       �                      @                                �|Y=@�t����?             A@        	                        ��*@����X�?             @       
                          �5@���Q��?             @        ������������������������       �                     �?                                  @@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                ���4@�>����?             ;@                                   @`2U0*��?             9@        ������������������������       �                      @                                �|�=@�nkK�?             7@                               ���@�8��8��?
             (@        ������������������������       �                     @                                  @@      �?              @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     &@                                `f&;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               .                    �?�?�'�@�?             C@              -                   �N@؇���X�?            �A@              ,                    �?�C��2(�?            �@@               %                  �>@H%u��?             9@        !       $                  Y>@���Q��?             @       "       #                 X��E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        &       +                   4W@P���Q�?             4@       '       (                  �oS@�����H�?             "@       ������������������������       �                     @        )       *                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        0       K                     �?�O��?�            �x@        1       J                    �?��
ц��?(            @P@       2       3                    �?�g�y��?&             O@        ������������������������       �        
             1@        4       I                 `f�D@�q�q�?            �F@       5       6                 03:@�g�y��?             ?@        ������������������������       �                     $@        7       F                 �T!@@����X�?             5@       8       E                   @>@������?             1@       9       B                 `fF<@�	j*D�?	             *@       :       A                   @L@z�G�z�?             $@       ;       <                 03k:@�����H�?             "@        ������������������������       �                     �?        =       >                   �C@      �?              @        ������������������������       �                     @        ?       @                   @G@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        C       D                   @K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        G       H                 �|�<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                     @        L       �                   �(@���/���?�            pt@       M       X                     @��W�'�?�            �l@        N       O                   �1@ �Cc}�?             <@        ������������������������       �                     �?        P       Q                    @�>����?             ;@        ������������������������       �                     @        R       W                    &@�����?             5@       S       V                    �?�KM�]�?	             3@        T       U                   �J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                      @        Y       n                    �?.p����?�            @i@        Z       [                 ��@���Q��?            �A@        ������������������������       �                      @        \       ]                    �?|��?���?             ;@        ������������������������       �                     @        ^       m                    �?���|���?             6@       _       d                 �?�@�z�G��?             4@        `       c                   �7@      �?              @        a       b                    4@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        e       j                    9@�q�q�?             (@       f       g                  �#@؇���X�?             @       ������������������������       �                     @        h       i                    4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        k       l                    A@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        o       �                   @@@ w���?i            �d@       p       �                 �?�@���� �?W             a@       q       �                 ��@`��F:u�?7            �U@       r       s                    7@�:�]��?            �I@        ������������������������       �                     .@        t                        �|Y=@�����H�?             B@        u       ~                    ;@�z�G��?             $@       v       w                    �?�<ݚ�?             "@        ������������������������       �                     �?        x       }                   �8@      �?              @       y       |                 `fF@���Q��?             @       z       {                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���@ ��WV�?             :@        ������������������������       �                     0@        ������������������������       �ףp=
�?             $@        ������������������������       �                     B@        �       �                 �|�=@���c�H�?             �H@       �       �                 ���"@�T|n�q�?            �E@       �       �                   �3@$G$n��?            �B@        �       �                 0S5 @����X�?             ,@        �       �                   �2@      �?              @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                    <@�nkK�?             7@        �       �                 pf� @�C��2(�?             &@       ������������������������       �                     "@        �       �                 @3�!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             (@        �       �                   �<@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 ��l!@�q�q�?             @       �       �                   �?@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     ?@        �       �                    �?@��Pl3�?:            @X@       �       �                 �|=@�G�z�?-             T@        �       �                    �?ףp=
�?             >@        �       �                     @���Q��?             @       �       �                    :@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @`2U0*��?             9@       ������������������������       �                     0@        �       �                 �T�C@�����H�?             "@       ������������������������       �                     @        �       �                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?z�):���?             I@        �       �                   �*@���7�?             6@       �       �                     @@4և���?             ,@       �       �                 ��Y)@�8��8��?             (@        ������������������������       �                      @        �       �                   �B@ףp=
�?             $@       ������������������������       �                      @        �       �                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                     @@4և���?             <@       �       �                   @A@P���Q�?             4@        �       �                    @@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �        	             *@        �       �                 0��A@      �?              @        ������������������������       �                     @        �       �                 �|�>@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    B@ҳ�wY;�?             1@       �       �                    �?�C��2(�?	             &@        ������������������������       �                     @        �       �                    �?r�q��?             @       �       �                     @z�G�z�?             @        ������������������������       �                      @        �       �                 `f7@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       >                   @�eH&b��?�            �m@       �       3                   @r�p���?�            �l@       �       �                    �?��>��?�            �i@        �       �                    �? s�n_Y�?#             J@       �       �                    �?Pa�	�?            �@@       �       �                   @0@ ��WV�?             :@        �       �                     @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     @        �       �                     �?�\��N��?             3@        �       �                 p"�X@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��3@�	j*D�?
             *@       �       �                    7@      �?              @        ������������������������       �                      @        �       �                 03�-@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �                          �?�@����?a            @c@       �       �                     @l�Ӑ���?2            �U@        �       �                    @��S�ۿ?            �F@        ������������������������       �                     �?        �       �                     �?���7�?             F@       ������������������������       �                     6@        �       �                    �?�C��2(�?             6@       �       �                    �?�KM�]�?	             3@        �       �                   �9@      �?              @        ������������������������       �                     @        �       �                   �7@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        �                          �?�D����?             E@       �       �                 P��%@��%��?            �B@        �       �                    4@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �                       �|�<@X�<ݚ�?             ;@        �       �                    �?      �?              @        ������������������������       �                     @        �                           @      �?             @       �       �                 P��)@�q�q�?             @        ������������������������       �                     �?        �                        ��/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                 @�����?             3@                             �|�=@      �?             0@        ������������������������       �                     @                                �@@X�<ݚ�?             "@                               �>@և���X�?             @        ������������������������       �                     �?        	      
                03C3@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                              �|Y?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �@@��y�:�?/            �P@                                �?�<ݚ�?             �F@                                 �?H%u��?             9@       ������������������������       �                     3@                              �|�<@      �?             @       ������������������������       �                     @        ������������������������       �                     @                              03�3@��Q��?             4@                                 +@      �?             $@       ������������������������       �                     @        ������������������������       �                     @                                 �?z�G�z�?             $@                                1@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        !      .                   �?�eP*L��?             6@       "      #                 x#J@      �?             2@        ������������������������       �                     @        $      +                   �?���Q��?	             .@       %      *                   F@�q�q�?             (@       &      '                `f�N@�����H�?             "@       ������������������������       �                     @        (      )                  �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ,      -               �G�A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        /      0                   &@      �?             @        ������������������������       �                      @        1      2                  �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        4      7                   �?�8��8��?             8@        5      6                   @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        8      =                   @@4և���?
             ,@       9      :                   �?�C��2(�?             &@       ������������������������       �                     "@        ;      <                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �*       h�h))��}�(h,h/h0M?KK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?����/��?��؊���?�������?333333�?�a�a�?��y��y�?      �?      �?              �?      �?        <<<<<<�?�?�m۶m��?�$I�$I�?333333�?�������?              �?      �?      �?      �?                      �?      �?        �Kh/��?h/�����?���Q��?{�G�z�?      �?        �Mozӛ�?d!Y�B�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?      �?              �?              �?      �?              �?      �?        y�5���?������?�$I�$I�?۶m۶m�?F]t�E�?]t�E�?���Q��?)\���(�?�������?333333�?      �?      �?              �?      �?              �?        �������?ffffff�?�q�q�?�q�q�?              �?      �?      �?              �?      �?                      �?              �?      �?                      �?����S��?����X�?�؉�؉�?�;�;�?��{���?�B!��?              �?UUUUUU�?UUUUUU�?�B!��?��{���?      �?        �$I�$I�?�m۶m��?�?xxxxxx�?;�;��?vb'vb'�?�������?�������?�q�q�?�q�q�?              �?      �?      �?              �?�������?�������?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?              �?                      �?�����?��a�Ϳ�?�|���?[�#P��?%I�$I��?۶m۶m�?              �?�Kh/��?h/�����?      �?        =��<���?�a�a�?�k(���?(�����?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �2|#
L�?:5r���?�������?333333�?              �?{	�%���?	�%����?              �?]t�E]�?F]t�E�?ffffff�?333333�?      �?      �?      �?      �?      �?                      �?      �?        �������?�������?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?                      �?W��1 �?E���w��?xxxxxx�?<<<<<<�?�u�7[��?Ȥx�L��?}}}}}}�?�?      �?        �q�q�?�q�q�?ffffff�?333333�?9��8���?�q�q�?      �?              �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?O��N���?;�;��?      �?        �������?�������?      �?        4և����?/�����?���)k��?6eMYS��?к����?���L�?�m۶m��?�$I�$I�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        �Mozӛ�?d!Y�B�?]t�E�?F]t�E�?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        ��4l7��?�n�'�i�?�������?�������?�������?�������?333333�?�������?      �?      �?      �?                      �?              �?���Q��?{�G�z�?      �?        �q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        H�z�G�?q=
ףp�?F]t�E�?�.�袋�?�$I�$I�?n۶m۶�?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?      �?      �?                      �?              �?              �?n۶m۶�?�$I�$I�?ffffff�?�������?۶m۶m�?�$I�$I�?      �?              �?      �?      �?              �?      �?      �?              �?      �?      �?                      �?�������?�������?F]t�E�?]t�E�?              �?UUUUUU�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?UUUUUU�?              �?      �?        �r�����?�F" >��?�%��~�?m5x�@�?����?�	����?;�;��?�;�;�?|���?|���?;�;��?O��N���?�������?�������?              �?      �?                      �?              �?y�5���?�5��P�?UUUUUU�?�������?              �?      �?        vb'vb'�?;�;��?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �Y�	qV�?S{���?/�I���?�7[�~��?�?�������?      �?        F]t�E�?�.�袋�?              �?F]t�E�?]t�E�?(�����?�k(���?      �?      �?              �?�������?333333�?      �?                      �?              �?              �?�0�0�?z��y���?���L�?}���g�?�������?�������?              �?      �?        �q�q�?r�q��?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        ^Cy�5�?Q^Cy��?      �?      �?              �?�q�q�?r�q��?�$I�$I�?۶m۶m�?      �?              �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �@��~�?~5&��?9��8���?�q�q�?)\���(�?���Q��?      �?              �?      �?      �?                      �?�������?ffffff�?      �?      �?              �?      �?        �������?�������?�m۶m��?�$I�$I�?              �?      �?              �?        ]t�E�?t�E]t�?      �?      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?        n۶m۶�?�$I�$I�?]t�E�?F]t�E�?      �?              �?      �?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ4�phG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM	hjh))��}�(h,h/h0M	��h2h3h4hph<�h=Kub������       z                     @�C�"���?�           8�@               ]                  x#J@��.k���?�            0t@                                  �?�R�Srq�?�            `m@               	                    �?P���Q�?/             T@                                    �?�����H�?             "@                                  �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        
                          �*@0z�(>��?'            �Q@                                   �?      �?             8@                                  �?R���Q�?             4@        ������������������������       �                     @                                `f�)@@�0�!��?
             1@                                 �J@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?                                   :@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �G@               N                    �?�����?]            `c@              /                 ��$:@�p ��?J            �^@                                  5@hA� �?,            �Q@                                  �2@z�G�z�?             @        ������������������������       �                     @                                  �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �)@��ɉ�?(            @P@        ������������������������       �                     6@        !       "                     �? �#�Ѵ�?            �E@        ������������������������       �                     @        #       $                 �|Y<@P���Q�?             D@        ������������������������       �                     .@        %       (                 �|�=@HP�s��?             9@        &       '                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        )       .                   �*@���7�?             6@       *       +                   @D@@4և���?	             ,@       ������������������������       �                     $@        ,       -                    G@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        0       9                    �?�#ʆA��?            �J@        1       8                  Y>@����X�?             ,@        2       7                 �|�=@�q�q�?             @       3       4                 �|�;@z�G�z�?             @        ������������������������       �                      @        5       6                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        :       I                   �F@�(�Tw��?            �C@       ;       H                   `@@�n_Y�K�?             :@       <       G                   @>@����X�?             ,@       =       D                 `fF<@���|���?             &@       >       ?                 03k:@      �?              @        ������������������������       �                      @        @       A                 �|�<@�q�q�?             @        ������������������������       �                     @        B       C                 X��B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        E       F                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        J       M                    J@$�q-�?	             *@        K       L                   �G@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        O       V                    :@      �?             @@       P       U                    �?b�2�tk�?
             2@       Q       R                    *@j���� �?	             1@        ������������������������       �                      @        S       T                    �?��S���?             .@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        W       X                    �?@4և���?	             ,@        ������������������������       �                     @        Y       Z                   �@@؇���X�?             @       ������������������������       �                     @        [       \                    0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ^       y                    @�~�4_��?8             V@       _       `                    �?�/,Tg�?6             U@       ������������������������       �                    �G@        a       x                   @I@��+��?            �B@       b       i                    �?����"�?             =@        c       d                 �|Y<@X�<ݚ�?             "@        ������������������������       �                     @        e       h                    �?r�q��?             @       f       g                 p�w@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        j       w                   �G@�z�G��?             4@       k       v                    �?���Q��?
             .@       l       u                    �?X�Cc�?	             ,@       m       n                    6@�n_Y�K�?             *@        ������������������������       �                      @        o       t                   �E@���!pc�?             &@       p       s                    >@�����H�?             "@        q       r                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        {       �                    �?�Ra�`��?�            @x@        |       �                    �?ד�w��?K            �^@        }       �                 X�,A@�p ��?            �D@       ~       �                    �?�˹�m��?             C@               �                    �?�θ�?	             *@       �       �                   �,@�q�q�?             "@        ������������������������       �                     @        �       �                 �%@���Q��?             @        ������������������������       �                     �?        �       �                   �7@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     9@        ������������������������       �                     @        �       �                    �?��]�T��?4            �T@       �       �                    @|��?���?%             K@        �       �                    �?؇���X�?             @        ������������������������       �                      @        �       �                     @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�=@�[�IJ�?             �G@       �       �                    �?      �?             D@       �       �                   �@�4�����?             ?@        �       �                    8@�z�G��?	             $@       �       �                   �2@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �9@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �)@؇���X�?             5@       ������������������������       �                     &@        �       �                    �?�z�G��?             $@       �       �                 03�0@և���X�?             @       �       �                 �|�;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �*@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��9$@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                     @      �?             @       �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �̼6@؇���X�?             <@        ������������������������       �                     @        �       �                 ��T?@`2U0*��?             9@       ������������������������       �                     1@        �       �                    @      �?              @        ������������������������       �                     @        �       �                 ���A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���[��?�            �p@       �       �                    �?8�ƨxt�?�            �k@       �       �                 �|Y=@��v����?s             i@        �       �                   �<@�~6�]�?4            @U@       �       �                    �?     ��?0             T@        �       �                    /@�q�q�?             .@        ������������������������       �                     @        �       �                   �7@r�q��?             (@        ������������������������       �                     "@        �       �                   �9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �:@$�q-�?+            @P@       �       �                   �3@h㱪��?&            �K@        �       �                   �1@�����H�?             2@        ������������������������       �                     @        �       �                 �?�@8�Z$���?
             *@        ������������������������       �                     @        �       �                   �2@�<ݚ�?             "@        �       �                 ��Y @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `�8"@؇���X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                    �B@        �       �                 �� @�z�G��?             $@        ������������������������       �                     @        �       �                   �;@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?,Z0R�??             ]@        ������������������������       �                     .@        �       �                   �@��T�u��?8            @Y@        �       �                    �?�T|n�q�?            �E@        �       �                 ���@      �?             0@        ������������������������       �                     @        ������������������������       �"pc�
�?             &@        �       �                 �&B@�+$�jP�?             ;@       �       �                 ��@�8��8��?             8@       ������������������������       �                     0@        �       �                 �|Y>@      �?              @        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    ?@XB���?!             M@       �       �                 ��) @ �#�Ѵ�?            �E@       ������������������������       �                    �A@        �       �                 pf� @      �?              @        ������������������������       �                     �?        �       �                    �?؇���X�?             @        ������������������������       �                     �?        �       �                 �|�=@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             .@        ������������������������       �                     4@        �                           @�zv�X�?             F@        �       �                    �?�t����?	             1@        �       �                 8#�2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                     @�θ�?             *@        ������������������������       �                     @        �       �                 ��T?@      �?             @       ������������������������       �                     @        ������������������������       �                     @                                  @�+$�jP�?             ;@                                �?X�Cc�?             ,@        ������������������������       �                     @                                 �?ףp=
�?             $@        ������������������������       �                     �?                                 )@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             *@        �*       h�h))��}�(h,h/h0M	KK��h2h3h4hVh<�h=Kub�������������[�e�?���I54�?�?�������?���R�?	��jZ��?�������?ffffff�?�q�q�?�q�q�?      �?      �?              �?      �?                      �?H���@��?�ԓ�ۥ�?      �?      �?333333�?333333�?              �?�������?ZZZZZZ�?F]t�E�?]t�E�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?���ۡ�?y�W�x�?Q��+Q�?��+Q��?���?_�_�?�������?�������?      �?              �?      �?              �?      �?        ?�?��? �����?      �?        �/����?�}A_Ч?      �?        ffffff�?�������?      �?        q=
ףp�?{�G�z�?UUUUUU�?UUUUUU�?      �?                      �?�.�袋�?F]t�E�?n۶m۶�?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        e�Cj���?5�x+��?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �o��o��?� � �?;�;��?ى�؉��?�$I�$I�?�m۶m��?F]t�E�?]t�E]�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �؉�؉�?;�;��?�������?UUUUUU�?      �?                      �?      �?              �?      �?�8��8��?9��8���?�������?ZZZZZZ�?      �?        �?�������?      �?                      �?      �?        n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        ��.���?]t�E�?=��<���?1�0��?              �?�S�n�?*�Y7�"�?�i��F�?	�=����?r�q��?�q�q�?              �?�������?UUUUUU�?�������?�������?      �?                      �?      �?        333333�?ffffff�?�������?333333�?�m۶m��?%I�$I��?ى�؉��?;�;��?      �?        t�E]t�?F]t�E�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?                      �?      �?                      �?_\����?BG����?.����-�?鰑��?��+Q��?Q��+Q�?^Cy�5�?��P^Cy�?�؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?              �?333333�?�������?              �?      �?      �?      �?                      �?              �?              �?      �?        KԮD�J�?jW�v%j�?{	�%���?	�%����?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?        ���
b�?m�w6�;�?      �?      �?���Zk��?��RJ)��?333333�?ffffff�?�$I�$I�?۶m۶m�?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?        ffffff�?333333�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?              �?        �q�q�?r�q��?              �?      �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?      �?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?              �?���Q��?{�G�z�?      �?              �?      �?      �?              �?      �?              �?      �?        �T�ѯ�?�ѯz�@�?�*�*�?�F�F�?5&����?*g��1�?999999�?�?      �?      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�؉�؉�?;�;��?־a���?��)A��?�q�q�?�q�q�?      �?        ;�;��?;�;��?      �?        9��8���?�q�q�?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?        ffffff�?333333�?      �?              �?      �?              �?      �?        �������?333333�?              �?      �?        �FX�i��?	�=��ܳ?      �?        Y�&�?:5r�϶?���)k��?6eMYS��?      �?      �?      �?        /�袋.�?F]t�E�?/�����?B{	�%��?UUUUUU�?UUUUUU�?      �?              �?      �?333333�?�������?      �?                      �?GX�i���?�{a���?�/����?�}A_Ч?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?      �?                      �?      �?              �?        ��.���?�袋.��?�������?�������?      �?      �?              �?      �?        �؉�؉�?ى�؉��?              �?      �?      �?      �?                      �?/�����?B{	�%��?%I�$I��?�m۶m��?              �?�������?�������?      �?        �q�q�?�q�q�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJLxhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM1hjh))��}�(h,h/h0M1��h2h3h4hph<�h=Kub������       h                    �?��l�Qf�?�           8�@               g                    @��"�y��?            �g@              $                   �9@�]$>��?~            �g@               #                    @~���L0�?            �H@                                  �?�q�q�?             H@                                 �1@�<ݚ�?             ;@        ������������������������       �                      @                                   5@�����?             3@        	       
                    �?�q�q�?             @        ������������������������       �                      @                                �{@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                   �?8�Z$���?             *@       ������������������������       �                     "@                                (SE&@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                �x"@�ՙ/�?             5@        ������������������������       �                      @                                 �U�X@�����?             3@                                    @r�q��?	             (@        ������������������������       �                     @                                �&�)@����X�?             @        ������������������������       �                     @                                   �?      �?             @                                  �?�q�q�?             @                                 �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        !       "                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        %       2                    �?&ޑ���?_            �a@        &       '                     @�1�`jg�?&            �K@       ������������������������       �                    �@@        (       /                    �?��2(&�?             6@       )       ,                 �YU&@�t����?             1@       *       +                    �?��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        -       .                 03�-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        0       1                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        3       J                 03�-@@�0�!��?9            @U@       4       A                    �?Hm_!'1�?            �H@       5       6                     @ 	��p�?             =@        ������������������������       �                      @        7       @                 �|�=@�>����?             ;@       8       ?                 ��� @�����H�?             2@       9       >                   @@"pc�
�?             &@       :       ;                 ���@ףp=
�?             $@        ������������������������       �                     @        <       =                 �|=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        B       I                 X��A@ףp=
�?             4@       C       D                  s�@�t����?
             1@        ������������������������       �                     @        E       H                    �?8�Z$���?             *@       F       G                 ��(@"pc�
�?             &@       ������������������������       ��<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        K       \                 �|�=@<ݚ)�?             B@        L       M                 ��.@      �?             4@        ������������������������       �                     @        N       O                 ��$1@      �?             0@        ������������������������       �                     @        P       Q                 03�7@��
ц��?	             *@        ������������������������       �                     @        R       U                 �|Y<@�z�G��?             $@        S       T                 Ъb@      �?             @        ������������������������       �                      @        ������������������������       �                      @        V       [                    �?r�q��?             @       W       X                 �ܵ<@z�G�z�?             @        ������������������������       �                      @        Y       Z                 03SA@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ]       f                    �?      �?             0@       ^       e                     �?ףp=
�?	             $@       _       `                    �?      �?              @       ������������������������       �                     @        a       b                   @G@�q�q�?             @        ������������������������       �                     �?        c       d                   �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        i                           �?V|�9�j�?D           @�@       j       �                    �?`S2(��?�            �x@        k       r                  �#@V��N��?9            �W@        l       m                 ���@8����?             7@        ������������������������       �                     @        n       o                   �9@z�G�z�?             4@       ������������������������       �                     (@        p       q                    ;@      �?              @        ������������������������       �                     @        ������������������������       �                     @        s       �                 `fF:@��UV�?+            �Q@       t       �                 03�1@z�G�z�?            �F@       u       �                     @<���D�?            �@@       v                          �*@؇���X�?             5@       w       z                    :@     ��?             0@        x       y                   �4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        {       ~                   �'@$�q-�?	             *@       |       }                   �J@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�8��8��?             (@        �       �                 �[$@z�G�z�?             @        ������������������������       �                      @        �       �                 ��&@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?             (@       �       �                     @�<ݚ�?             "@       �       �                  ��9@      �?              @        ������������������������       �                     �?        �       �                    �?؇���X�?             @        ������������������������       �                     �?        �       �                   �E@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        �       �                     �?,:#\��?�            �r@        �       �                    �?��>4և�?#             L@       �       �                    �?��}*_��?"             K@       �       �                   �9@�n_Y�K�?            �C@        ������������������������       �                      @        �       �                    D@�g�y��?             ?@        �       �                 X�,@@�	j*D�?             *@       �       �                 �|Y=@���|���?             &@       �       �                   �<@      �?             @       �       �                 `f�D@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `fF<@����X�?             @        ������������������������       �                     �?        �       �                 @�x_@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �G@�q�q�?             2@        ������������������������       �                     @        �       �                   �J@�eP*L��?	             &@        ������������������������       �                     @        �       �                  )?@����X�?             @        �       �                    R@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �B@�q�q�?             .@        ������������������������       �                     @        �       �                 0�nL@      �?             $@        ������������������������       �                     @        �       �                 03�U@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�R����?�            @n@       �       �                     @�j��b�?�            �m@        �       �                   @A@$Q�q�?$            �O@       �       �                    �?dP-���?            �G@       �       �                    @@�KM�]�?             C@       �       �                   �3@ >�֕�?            �A@       �       �                    5@��S�ۿ?             >@        �       �                    &@�����H�?             "@        ������������������������       �z�G�z�?             @        ������������������������       �                     @        �       �                 �|�<@���N8�?             5@        ������������������������       �                     (@        �       �                   �'@�����H�?             "@       ������������������������       �                     @        �       �                 �|�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �        
             0@        �       �                    �?��㨇,�?q            �e@       �       �                 �T�C@|�@�E-�?i             d@       �       �                 @3�@�f���?g            �c@       �       �                   �?@�=C|F�?8            �U@       �       �                   �7@      �?*             P@        ������������������������       �                     6@        �       �                 ���@�����?             E@        �       �                   �8@      �?             @        �       �                 �&b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y=@������?             B@        ������������������������       �        
             1@        �       �                  sW@�}�+r��?             3@        �       �                 �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        �       �                 �Y5@8����?             7@       ������������������������       �                     (@        �       �                   �@���|���?             &@        ������������������������       �                     �?        �       �                 �?�@���Q��?             $@        ������������������������       �                     �?        �       �                   �A@�q�q�?             "@       ������������������������       �      �?             @        ������������������������       �                     @        �       �                 pf!@hA� �?/            �Q@        ������������������������       �                    �A@        �       �                 ���!@�#-���?            �A@        �       �                    8@����X�?             @        ������������������������       �                     @        �       �                 �|Y<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 `�X#@h�����?             <@       �       �                   �=@�IєX�?             1@       ������������������������       �        	             (@        �       �                   �?@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                 �|�>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    5@      �?             (@        �       �                  s�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                              03s;@     ��?O             `@                                �;@`�Q��?!             I@                               �2@��� ��?             ?@                                -@�㙢�c�?             7@             
                   @      �?             0@                                 @      �?              @       ������������������������       �                     @              	                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                 �?����X�?             @                                �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @                                 �?p�ݯ��?             3@                                �?      �?	             0@                                 @X�<ݚ�?             "@        ������������������������       �                     �?                              `fv1@      �?              @        ������������������������       �                     @                                  @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @              *                    @�	j*D�?.            �S@              )                  �J@     ��?             @@             "                   @H%u��?             9@               !                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        #      (                   �?���}<S�?             7@        $      %                  �B@z�G�z�?             $@       ������������������������       �                     @        &      '                  @D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             *@        ������������������������       �                     @        +      ,                   @�nkK�?             G@        ������������������������       �                     .@        -      0                ���A@`Jj��?             ?@        .      /                ��T?@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     4@        �*       h�h))��}�(h,h/h0M1KK��h2h3h4hVh<�h=Kub������������}<����?�/���?o��2�|�?H���A�?��!s���?�oF��?������?����>4�?�������?�������?�q�q�?9��8���?              �?^Cy�5�?Q^Cy��?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?;�;��?;�;��?              �?      �?      �?              �?      �?        �a�a�?�<��<��?      �?        ^Cy�5�?Q^Cy��?UUUUUU�?�������?              �?�$I�$I�?�m۶m��?              �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?              �?        �������?���?�־a�?A��)A�?              �?t�E]t�?��.���?�?<<<<<<�?�?�������?              �?      �?              �?      �?      �?                      �?�������?�������?      �?                      �?ZZZZZZ�?�������?Y�Cc�?9/���?������?�{a���?      �?        �Kh/��?h/�����?�q�q�?�q�q�?/�袋.�?F]t�E�?�������?�������?      �?        �������?�������?      �?              �?      �?              �?      �?              �?        �������?�������?<<<<<<�?�?      �?        ;�;��?;�;��?/�袋.�?F]t�E�?9��8���?�q�q�?      �?              �?              �?        ��8��8�?�8��8��?      �?      �?              �?      �?      �?      �?        �;�;�?�؉�؉�?              �?ffffff�?333333�?      �?      �?              �?      �?        �������?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?                      �?��Z��Z�?��J��J�?������?�>4և��?��
br�?����F}�?d!Y�B�?8��Moz�?              �?�������?�������?      �?              �?      �?              �?      �?        6��9�?2~�ԓ��?�������?�������?|���?|���?�$I�$I�?۶m۶m�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?�؉�؉�?�$I�$I�?۶m۶m�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?�q�q�?9��8���?      �?      �?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?              �?      �?              �?              �?                      �?���v�?�t�%��?۶m۶m�?I�$I�$�?_B{	�%�?B{	�%��?;�;��?ى�؉��?      �?        �B!��?��{���?;�;��?vb'vb'�?F]t�E�?]t�E]�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?        ]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?�m۶m��?�$I�$I�?      �?                      �?              �?�������?���!pc�?�N��?��/���?~��}���?AA�?�����F�?W�+�ɵ?�k(���?(�����?��+��+�?�A�A�?�������?�?�q�q�?�q�q�?�������?�������?      �?        ��y��y�?�a�a�?      �?        �q�q�?�q�q�?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?              �?        ۜ��L�?�'�j��?�O���?���G��?̟�Ѐ%�?�Kz�Ӷ?�C��:��?J��/�?      �?      �?      �?        =��<���?�a�a�?      �?      �?      �?      �?      �?                      �?      �?        �q�q�?�q�q�?      �?        �5��P�?(�����?      �?      �?              �?      �?              �?        d!Y�B�?8��Moz�?      �?        F]t�E�?]t�E]�?              �?�������?333333�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?���?_�_�?      �?        �A�A�?_�_�?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?        �m۶m��?�$I�$I�?�?�?      �?        �������?�������?              �?      �?              �?              �?      �?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?              �?             ��?      �?{�G�z�?��(\���?�B!��?�{����?d!Y�B�?�7��Mo�?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?�m۶m��?�������?333333�?              �?      �?                      �?              �?^Cy�5�?Cy�5��?      �?      �?r�q��?�q�q�?              �?      �?      �?      �?        �������?333333�?              �?      �?              �?                      �?vb'vb'�?;�;��?      �?      �?���Q��?)\���(�?      �?      �?              �?      �?        d!Y�B�?ӛ���7�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �Mozӛ�?d!Y�B�?      �?        ���{��?�B!��?/�袋.�?F]t�E�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW��8hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       d                    �?H���I�?�           8�@               !                     @���N8�?�            �o@                                  �?�X�<ݺ?U             b@                                  L@��S�ۿ?9            @Z@              
                   �;@p�qG�?5             X@               	                   �7@ܷ��?��?             =@                                   )@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     3@                                   �?0�,���?$            �P@                                  �? 7���B�?             K@                                  �F@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?                                   -@ qP��B�?            �E@                               `f�)@(;L]n�?             >@        ������������������������       �                     (@                                  �B@�X�<ݺ?             2@       ������������������������       �                     0@                                   D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �        	             *@                                  �L@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @                                ���a@ ���J��?            �C@       ������������������������       �                     ?@                                    !@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        "       Q                    �?|��?���?E             [@       #       4                    �?^�JB=�?3            @T@        $       +                   �2@b�h�d.�?            �A@        %       &                    �?�q�q�?             "@        ������������������������       �                     @        '       *                 `�@1@      �?             @       (       )                 P��+@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ,       /                    �?ȵHPS!�?             :@        -       .                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        0       3                    �?�C��2(�?             6@       1       2                 ���@      �?             0@        ������������������������       �                      @        ������������������������       �        
             ,@        ������������������������       �                     @        5       P                    �?(옄��?             G@       6       ;                    3@�p ��?            �D@        7       :                 ��!@      �?              @        8       9                 P��@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        <       A                 P�@4���C�?            �@@        =       @                 ��@�n_Y�K�?             *@       >       ?                 �|Y:@�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        B       I                    �?�z�G��?             4@       C       D                   �9@����X�?	             ,@       ������������������������       �                     "@        E       F                    �?z�G�z�?             @        ������������������������       �                     �?        G       H                 `f�/@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        J       K                   �&@�q�q�?             @        ������������������������       �                      @        L       M                    �?      �?             @        ������������������������       �                     �?        N       O                 `fV6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        R       U                    �?�<ݚ�?             ;@        S       T                 �|�:@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        V       Y                    �?�d�����?             3@        W       X                 `f7@      �?             @        ������������������������       �                     @        ������������������������       �                     @        Z       [                    @8�Z$���?             *@        ������������������������       �                     @        \       ]                 ���3@����X�?             @        ������������������������       �                     �?        ^       c                 pf�C@r�q��?             @       _       `                    @�q�q�?             @        ������������������������       �                     �?        a       b                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        e       �                    �?��`��?           �|@       f       g                    $@�ɮ����?�            �v@        ������������������������       �                     @        h       �                     �?�:�^���?�            �v@        i       �                    @@2%ޑ��?'            �Q@       j       y                 ���=@      �?             B@       k       l                   �9@r�q��?             >@        ������������������������       �                     (@        m       x                    B@�E��ӭ�?             2@       n       w                 ���<@      �?             $@       o       v                 ��";@      �?              @       p       q                 03k:@���Q��?             @        ������������������������       �                     �?        r       s                    �?      �?             @        ������������������������       �                     �?        t       u                 �|�<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        z       {                    <@�q�q�?             @        ������������������������       �                     �?        |       �                  �>@���Q��?             @       }       ~                    �?      �?             @        ������������������������       �                     �?               �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��UO@�IєX�?             A@       ������������������������       �        
             3@        �       �                    �?�r����?             .@       �       �                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �       �                   @@@DK{22�?�             r@       �       �                 ��q1@����X��?�             l@       �       �                    �?�n���?�             k@        �       �                   �6@д>��C�?             =@        ������������������������       �                      @        �       �                 ���@�����H�?             ;@        ������������������������       �                     *@        �       �                 �|�=@d}h���?             ,@       �       �                   @@      �?             (@       ������������������������       �և���X�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@a��_�?r            `g@       �       �                   �<@���J��?<            �Y@        ������������������������       �                    �H@        �       �                     @�&=�w��?!            �J@        ������������������������       �                     &@        �       �                 �|Y=@���N8�?             E@        �       �                   @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�(\����?             D@        �       �                  s�@      �?             0@        ������������������������       �                     @        �       �                 ��(@�C��2(�?	             &@       ������������������������       �ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     8@        �       �                    �?��O���?6            @U@        ������������������������       �                     �?        �       �                     @�����?5             U@        �       �                    5@���}<S�?             7@        �       �                    &@�q�q�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �        	             1@        �       �                 ���#@\#r��?(            �N@       �       �                   �<@�����H�?$             K@        �       �                    1@�nkK�?             7@        �       �                 pFD!@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     3@        �       �                 ��) @�חF�P�?             ?@       �       �                 @3�@���7�?             6@        �       �                   �?@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             1@        �       �                 ��y @X�<ݚ�?             "@        ������������������������       �                      @        �       �                 �|Y=@����X�?             @        ������������������������       �                     �?        �       �                 �|�=@r�q��?             @        ������������������������       �                     @        �       �                 ���!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @        �       �                   �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     @���Q��?             @        ������������������������       �                     �?        �       �                    ;@      �?             @        ������������������������       �                      @        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @Pa�	�?(            �P@        �       �                    �?      �?             0@        ������������������������       �                      @        �       �                    �?@4և���?	             ,@       �       �                   @F@$�q-�?             *@        �       �                   �C@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?p���?             I@       �       �                 �?�@@��8��?             H@       ������������������������       �                     >@        �       �                   @D@�X�<ݺ?             2@       �       �                   @B@�����H�?             "@       ������������������������       �                     @        �       �                 ��	0@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        �       �                     �?�ț��*�?@            �W@        �       �                    �?      �?             6@       �       �                     @      �?             2@       �       �                 Ј�U@     ��?             0@       �       �                    �?�eP*L��?             &@        ������������������������       �                     @        �       �                    A@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �5@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���[@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �                         �C@z�z�7��?2            @R@       �                          �?Z���c��?*            �O@        �       �                    �?�����?             5@        ������������������������       �                     @        �       �                    �?�����H�?             2@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          �?@4և���?             ,@       �       �                     @�8��8��?	             (@        ������������������������       �                     @                                  5@؇���X�?             @                              �Y�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                 @0,Tg��?             E@                                 �?d}h���?	             ,@        ������������������������       �                      @        	      
                   �?�8��8��?             (@        ������������������������       �                     @                                 @z�G�z�?             @                              ���7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@        ������������������������       �                     $@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������Q�Ȟ���?^-n����?��y��y�?�a�a�?�q�q�?��8��8�?�?�������?�������?UUUUUU�?a���{�?��=���?333333�?ffffff�?              �?      �?                      �?g��1��?Ez�rv�?h/�����?	�%����?F]t�E�?]t�E�?              �?      �?        �}A_З?��}A�?�?�������?              �?�q�q�?��8��8�?              �?      �?      �?      �?                      �?              �?              �?�q�q�?9��8���?      �?                      �?�A�A�?��-��-�?              �?      �?      �?      �?                      �?	�%����?{	�%���?�2�tk~�?��E���?_�_��?;��:���?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?              �?      �?                      �?�؉�؉�?��N��N�?      �?      �?      �?                      �?F]t�E�?]t�E�?      �?      �?      �?                      �?              �?���,d�?ӛ���7�?8��18�?dp>�c�?      �?      �?      �?      �?              �?      �?                      �?m��&�l�?'�l��&�?ى�؉��?;�;��?]t�E�?t�E]t�?              �?      �?                      �?ffffff�?333333�?�m۶m��?�$I�$I�?      �?        �������?�������?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        9��8���?�q�q�?      �?      �?              �?      �?        Cy�5��?y�5���?      �?      �?              �?      �?        ;�;��?;�;��?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?        |&�{&��?f�f��?]��\���?�Q�Q�?              �?}�'}�'�?l�l��?�������?�A�A�?      �?      �?�������?UUUUUU�?      �?        �q�q�?r�q��?      �?      �?      �?      �?�������?333333�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?              �?�������?333333�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�?�?      �?        �������?�?UUUUUU�?UUUUUU�?              �?      �?              �?        ���Dɮ�?^�(ٵ��?�$I�$I�?n۶m۶�?r�q��?r�qǱ?a���{�?|a���?              �?�q�q�?�q�q�?      �?        I�$I�$�?۶m۶m�?      �?      �?�$I�$I�?۶m۶m�?      �?              �?        J����I�?a�2a�?______�?�?      �?        tHM0���?�x+�R�?      �?        ��y��y�?�a�a�?      �?      �?              �?      �?        333333�?�������?      �?      �?      �?        ]t�E�?F]t�E�?�������?�������?      �?              �?        �������?�?      �?        =��<���?�a�a�?ӛ���7�?d!Y�B�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        ��:��?XG��).�?�q�q�?�q�q�?�Mozӛ�?d!Y�B�?      �?      �?      �?      �?      �?              �?        �Zk����?��RJ)��?�.�袋�?F]t�E�?�������?�������?              �?      �?              �?        r�q��?�q�q�?              �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?      �?              �?      �?              �?      �?      �?      �?                      �?|���?|���?      �?      �?      �?        n۶m۶�?�$I�$I�?�؉�؉�?;�;��?�������?�������?      �?              �?      �?      �?              �?        \���(\�?{�G�z�?UUUUUU�?UUUUUU�?      �?        ��8��8�?�q�q�?�q�q�?�q�q�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?              �?        �~�-q��?�a�+�?      �?      �?      �?      �?      �?      �?t�E]t�?]t�E�?              �?      �?      �?              �?      �?        �������?�������?      �?                      �?      �?              �?      �?      �?                      �?ҤI�&M�?�lٲe��?Y�eY�e�?��i��i�?=��<���?�a�a�?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?        �y��y��?1�0��?۶m۶m�?I�$I�$�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?      �?                      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��UhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       b                    �?e�L��?�           8�@                                  �2@��,?S�?�            @n@                                    @F�����?            �F@                                ��Z@      �?	             0@       ������������������������       �                     *@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        	                           @l��[B��?             =@       
                        `f7@�q�q�?             8@                                �2@�z�G��?             4@                                  �?��
ц��?
             *@                                  �?�q�q�?	             (@                                  1@և���X�?             @       ������������������������       �                     @                                P��@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?���Q��?             @                                   &@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               a                    @���mf�?~            �h@              P                   @D@��_I(�?{            �g@              O                 ���7@�"ZN��?b            �b@              &                 �̌@:���u��?8            @S@                !                    8@H%u��?             9@        ������������������������       �                     &@        "       #                 ���@d}h���?	             ,@        ������������������������       �                      @        $       %                    �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        '       6                     @�	j*D�?*             J@        (       3                   `2@�㙢�c�?             7@       )       0                   �B@ףp=
�?             4@       *       /                   �9@�X�<ݺ?             2@        +       .                    �?�q�q�?             @       ,       -                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        1       2                   �,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        4       5                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        7       <                    �?�f7�z�?             =@        8       9                 �|Y=@ףp=
�?             $@        ������������������������       �                     @        :       ;                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        =       D                   �&@D�n�3�?             3@        >       C                 pf� @z�G�z�?             $@        ?       @                   �8@���Q��?             @        ������������������������       �                      @        A       B                 �?�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        E       J                 03�1@�q�q�?             "@       F       G                    �?r�q��?             @       ������������������������       �                     @        H       I                   �;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        K       L                 03C3@�q�q�?             @        ������������������������       �                     �?        M       N                 ���5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        *            �Q@        Q       `                     @�lg����?            �E@       R       _                 �DD@"pc�
�?            �@@        S       ^                    �?���Q��?
             .@       T       U                   @F@      �?             (@        ������������������������       �                     @        V       W                    �?�q�q�?             "@        ������������������������       �                      @        X       Y                     �?؇���X�?             @        ������������������������       �                      @        Z       ]                    (@z�G�z�?             @       [       \                   �J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     $@        ������������������������       �                     @        c       �                    �?�Y����?0           P}@        d       �                    �?��j���?0            �T@       e       �                 p�w@�����?#            �L@       f       k                   @@�E��ӭ�?"             K@        g       h                 03S@      �?             0@        ������������������������       �                     �?        i       j                   �6@�r����?             .@        ������������������������       �                      @        ������������������������       �        	             *@        l       m                 �� @P����?             C@        ������������������������       �                     @        n                            �?����X�?            �A@       o       p                 ��";@�c�Α�?             =@        ������������������������       �                     @        q       ~                    �?���B���?             :@       r       s                 ���=@�q�q�?             8@        ������������������������       �                      @        t       }                   �F@     ��?
             0@       u       |                    �?      �?              @       v       {                 `f�A@և���X�?             @       w       z                 X�lA@z�G�z�?             @       x       y                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                 �|�;@z�G�z�?             @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��
ц��?             :@       �       �                     �?�q�����?             9@        �       �                   �5@r�q��?             (@        ������������������������       �                     �?        �       �                   �H@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                     @8�Z$���?             *@       ������������������������       �                     "@        �       �                 03�-@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?Z�ڤ��?             x@        �       �                 X��A@�חF�P�?             ?@       �       �                  ��@z�G�z�?             9@        ������������������������       �                     @        �       �                    2@      �?             4@        ������������������������       �                     @        �       �                 03�7@     ��?             0@       �       �                 �|Y=@�q�q�?             .@        ������������������������       �                      @        �       �                   `3@�θ�?             *@       �       �                 ��(@r�q��?             (@       �       �                    �?�<ݚ�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��$:@�
d�<u�?�            0v@       �       �                    )@�c:��?�            @q@        ������������������������       �                     @        �       �                     @�X�<ݺ?�            �p@        �       �                     �?@�j;��?0            �Q@        ������������������������       �                     .@        �       �                    4@ �Cc}�?(             L@        �       �                    &@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                   @D@=QcG��?"            �G@       �       �                    �?�g�y��?             ?@       �       �                   �(@(;L]n�?             >@        ������������������������       �        
             ,@        �       �                    1@      �?             0@       �       �                 �|Y<@ףp=
�?             $@       ������������������������       �                     @        �       �                 �|�?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?
             0@       �       �                    F@؇���X�?             ,@        ������������������������       �      �?             @        ������������������������       �                     $@        ������������������������       �                      @        �       �                 `�X#@�����?~            �h@       �       �                    �?�}�+r��?k            `e@       �       �                   �?@�<� w�?c            �c@       �       �                 ���"@H�̱���?I            @_@       �       �                 �?$@ @|���?F            �^@        �       �                    7@������?            �B@       ������������������������       �                     2@        �       �                   �8@���y4F�?	             3@        ������������������������       �                     �?        �       �                 pf�@r�q��?             2@       ������������������������       �                     ,@        ������������������������       �      �?             @        �       �                 �?�@@�)�n�?1            @U@        ������������������������       �                    �D@        �       �                   �>@t��ճC�?             F@       �       �                   � @ �#�Ѵ�?            �E@       �       �                   �2@(;L]n�?             >@        �       �                    1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        �       �                 @�!@$�q-�?	             *@       �       �                   �7@؇���X�?             @       ������������������������       �                     @        �       �                 �|Y<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    =@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     A@        �       �                    �?�8��8��?             (@       �       �                 P�@�C��2(�?             &@       ������������������������       �                     @        �       �                    7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     <@        �                           �?H���I�?4            �S@       �       �                    @@П[;U��?%             M@        �       �                   �J@�����?             3@       �       �                 �|�<@؇���X�?	             ,@        ������������������������       �                     @        �       �                 `fF<@z�G�z�?             $@       �       �                 03k:@����X�?             @        ������������������������       �                     �?        �       �                    H@�q�q�?             @       �       �                 X��B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �Q@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �                         �;@�q�q�?            �C@        �                           �?      �?              @        �       �                    7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                              �|Y>@��a�n`�?             ?@        ������������������������       �                     "@                                �E@�X����?             6@                               x#J@      �?              @        ������������������������       �                      @        ������������������������       �                     @              	                ��#[@@4և���?
             ,@       ������������������������       �                     (@        
                        �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              ��T?@�����?             5@        ������������������������       �                     @                                 ;@�r����?
             .@                                5@�<ݚ�?             "@                                @      �?              @                                  @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������v�S(��?��X��?����|��?�ˠT�?؂-؂-�?�>�>��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ���=��?GX�i���?�������?�������?333333�?ffffff�?�؉�؉�?�;�;�?�������?�������?۶m۶m�?�$I�$I�?              �?      �?      �?              �?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?              �?        �H(m���?���W�?G��y�t�?��!�"�?�S�n�?E>�S��?qV~B���?dj`��?���Q��?)\���(�?              �?۶m۶m�?I�$I�$�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ;�;��?vb'vb'�?d!Y�B�?�7��Mo�?�������?�������?�q�q�?��8��8�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        a���{�?O#,�4��?�������?�������?              �?UUUUUU�?�������?              �?      �?        l(�����?(������?�������?�������?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�}A_��?}A_��?F]t�E�?/�袋.�?�������?333333�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?      �?              �?        ��¯�D�?���@���?�e�@	o�?o4u~�!�?Q^Cy��?^Cy�5�?�q�q�?r�q��?      �?      �?      �?        �������?�?              �?      �?        �P^Cy�?Q^Cy��?              �?�m۶m��?�$I�$I�?5�rO#,�?�{a���?              �?��؉���?ى�؉��?UUUUUU�?�������?      �?              �?      �?      �?      �?۶m۶m�?�$I�$I�?�������?�������?      �?      �?              �?      �?                      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?      �?                      �?              �?�;�;�?�؉�؉�?�p=
ף�?���Q��?UUUUUU�?�������?      �?        F]t�E�?]t�E�?              �?      �?        ;�;��?;�;��?      �?              �?      �?      �?                      �?      �?        ���
���?n����?�Zk����?��RJ)��?�������?�������?      �?              �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?ى�؉��?�؉�؉�?�������?UUUUUU�?9��8���?�q�q�?      �?      �?      �?              �?                      �?      �?              �?        B�E��?���3��?Y�B���?8��Moz�?              �?��8��8�?�q�q�?w�'�K�?H���@��?      �?        %I�$I��?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?        x6�;��?AL� &W�?��{���?�B!��?�������?�?      �?              �?      �?�������?�������?      �?              �?      �?              �?      �?              �?              �?              �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?              �?        Ym�큍�?t*) �'�?�5��P�?(�����?���c�?��N�©?�ʡE���?����Mb�?"XG��)�?�}�K�`�?��g�`��?к����?      �?        6��P^C�?(������?              �?�������?UUUUUU�?      �?              �?      �?�������?�?      �?        �E]t��?t�E]t�?�/����?�}A_Ч?�������?�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �؉�؉�?;�;��?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?]t�E�?F]t�E�?      �?              �?      �?              �?      �?              �?              �?        Q�Ȟ���?^-n����?�{a���?��=���?^Cy�5�?Q^Cy��?�$I�$I�?۶m۶m�?              �?�������?�������?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?              �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�c�1��?�s�9��?      �?        �E]t��?]t�E]�?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?      �?              �?      �?              �?      �?        =��<���?�a�a�?      �?        �������?�?9��8���?�q�q�?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��DphG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       b                    �?@t]q�V�?�           8�@               ]                    @��	�3��?�             m@              >                 �|�=@Ƶ�pD�?�             k@                                   @�����?X            �`@                                   �?�h����?%             L@        ������������������������       �        	             ,@                                   �?@4և���?             E@                                  �;@�r����?             .@       	       
                    �?      �?              @       ������������������������       �                     @                                  �9@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                   �? 7���B�?             ;@       ������������������������       �        
             .@                                   @�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@                                   �?�):u��?3            @S@                                   �?V������?            �B@                                  �?д>��C�?             =@                                   �?      �?             $@        ������������������������       �                     @                                �&�)@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@                                `�@1@      �?              @       ������������������������       �                     @        ������������������������       �                      @                1                    �?      �?             D@       !       ,                    �?      �?             8@       "       '                   �5@j���� �?             1@        #       $                    '@      �?              @        ������������������������       �                     @        %       &                 ���@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        (       +                   �@�����H�?             "@        )       *                 P��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        -       0                    ,@����X�?             @       .       /                    @      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        2       3                 P�@     ��?             0@        ������������������������       �                     �?        4       =                    �?�r����?             .@       5       <                 03�0@8�Z$���?	             *@       6       9                    �?      �?              @       7       8                 �|�;@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        :       ;                    -@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ?       R                    �?؇���X�?5             U@       @       A                   @B@�GN�z�?             F@        ������������������������       �                     4@        B       E                   �C@�q�q�?             8@        C       D                     �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        F       Q                    @������?             1@       G       N                 0#R;@     ��?             0@       H       I                     �?ףp=
�?             $@        ������������������������       �                      @        J       M                   �'@      �?              @        K       L                   �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        O       P                 ,w�U@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        S       \                    @P���Q�?             D@       T       [                    �? ���J��?            �C@       U       V                    @������?             B@       ������������������������       �                    �@@        W       Z                    @�q�q�?             @       X       Y                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ^       _                   �3@     ��?
             0@        ������������������������       �                     @        `       a                      @X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        c       �                     �?(a��0�?-           �}@        d       �                    �?     ��?<             X@       e       �                   @J@��}*_��?3            @T@       f       s                  �>@T�iA�?+            �Q@        g       h                 ��<:@��X��?             <@        ������������������������       �                     @        i       r                 �ܵ<@��2(&�?             6@       j       q                 ��";@z�G�z�?             .@       k       l                    �?$�q-�?             *@        ������������������������       �                      @        m       p                   @G@�C��2(�?             &@       n       o                   �C@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        t       �                    H@���N8�?             E@       u       ~                    �?�t����?             A@        v       }                    �?�q�q�?             "@       w       |                 X�lA@      �?              @       x       {                  �}S@r�q��?             @        y       z                 �|Y<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?               �                 03�U@`2U0*��?             9@       ������������������������       �                     2@        �       �                   �D@؇���X�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @       �       �                   �H@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�C��2(�?             &@        ������������������������       �                     �?        �       �                    R@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?z�G�z�?	             .@       �       �                   �7@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    =@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �                          �?H,Z�"��?�            �w@       �       �                     @H�/�.K�?�            �u@        �       �                    #@�<p���?8            �T@        ������������������������       �                     @        �       �                    �?p�|�i�?5             S@        ������������������������       �                     @        �       �                    �?hA� �?0            �Q@       �       �                   �*@�1�`jg�?'            �K@       �       �                    @��S�ۿ?             �F@        ������������������������       �                     @        �       �                    &@��(\���?             D@        �       �                   �5@ףp=
�?             $@        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                 `fF)@��S�ۿ?             >@        ������������������������       �                     @        �       �                 �|Y<@�8��8��?             8@        ������������������������       �                     $@        �       �                 �|�=@؇���X�?
             ,@        ������������������������       �                     �?        �       �                   @D@$�q-�?	             *@        ������������������������       �                     @        �       �                   �F@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        	             .@        �       �                    �?�$�^��?�            �p@       �       �                   �<@�n%����?�            �m@        �       �                 �?�@b �57�?D            �Y@       �       �                 �Y�@���J��?#            �I@        �       �                 ���@$�q-�?	             *@       ������������������������       �                     $@        �       �                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     C@        �       �                    �?ȵHPS!�?!             J@        ������������������������       �                     �?        �       �                   �2@�t����?             �I@        �       �                   �1@�z�G��?             $@       �       �                 pf� @      �?              @        ������������������������       �      �?             @        ������������������������       �                     @        �       �                 ��Y @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��p\�?            �D@       �       �                   �;@�7��?            �C@       �       �                   �:@�>����?             ;@       �       �                 0S5 @ ��WV�?             :@        �       �                    4@�C��2(�?             &@        ������������������������       �      �?              @        ������������������������       �                     "@        ������������������������       �        	             .@        ������������������������       �                     �?        ������������������������       �                     (@        �       �                 pf(@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���>���?R            �`@       �       �                 �|Y=@t�7��?M             _@        ������������������������       �                     @        �       �                  s�@�ݜ�?J            @]@        �       �                 ���@��Y��]�?            �D@       ������������������������       �                     <@        �       �                 �|�=@$�q-�?             *@       �       �                    �?�8��8��?             (@        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @@@>A�F<�?3             S@       �       �                   �>@x��}�?"            �K@       �       �                    �?*
;&���?             G@        ������������������������       �                     @        �       �                  sW@r�q��?             E@        �       �                 ��@և���X�?             ,@       ������������������������       �����X�?             @        ������������������������       �և���X�?             @        �       �                 ��)"@h�����?             <@       ������������������������       �                     7@        �       �                    (@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �&B@�q�q�?             "@        ������������������������       �                     �?        �       �                 P�@      �?              @        ������������������������       �                     �?        �       �                   �?@����X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        �       �                    �?���N8�?             5@        ������������������������       �                     @        �       �                   @C@�IєX�?             1@       ������������������������       �                     (@        �       �                 @3�@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    )@     ��?             @@        ������������������������       �                     @        �                       �|�?@8�Z$���?             :@        �                           3@�	j*D�?             *@       ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     *@                                 @      �?             @@                                 �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ;@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������
���?�;����?�=���?<ọ'|�?�Tx*<�?��a��z�?E,�T��?�iu�՝�?۶m۶m�?�$I�$I�?              �?�$I�$I�?n۶m۶�?�?�������?      �?      �?              �?      �?      �?              �?      �?                      �?h/�����?	�%����?              �?UUUUUU�?UUUUUU�?      �?                      �?5�wL��?�'�Y�	�?o0E>��?�g�`�|�?|a���?a���{�?      �?      �?              �?�������?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?      �?      �?      �?      �?�������?ZZZZZZ�?      �?      �?              �?�������?333333�?              �?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?      �?              �?�������?�?;�;��?;�;��?      �?      �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �$I�$I�?۶m۶m�?]t�E�?�袋.��?              �?�������?�������?۶m۶m�?�$I�$I�?              �?      �?        �?xxxxxx�?      �?      �?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?ffffff�?�A�A�?��-��-�?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?      �?              �?      �?      �?        �q�q�?r�q��?              �?      �?        �&䅭��?�eo�I��?      �?      �?_B{	�%�?B{	�%��?�+��+��?;��:���?%I�$I��?n۶m۶�?      �?        t�E]t�?��.���?�������?�������?;�;��?�؉�؉�?              �?F]t�E�?]t�E�?�������?�������?              �?      �?                      �?      �?                      �?�a�a�?��y��y�?<<<<<<�?�?UUUUUU�?UUUUUU�?      �?      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        ���Q��?{�G�z�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?]t�E�?F]t�E�?      �?        �������?�������?      �?                      �?�������?�������?�������?�������?              �?      �?        333333�?�������?              �?      �?        z�t�1��?�-�9k�?/ 6����?E'���?}���|�?�����?              �?�k(����?^Cy�5�?      �?        ���?_�_�?A��)A�?�־a�?�������?�?      �?        �������?333333�?�������?�������?UUUUUU�?UUUUUU�?      �?        �������?�?      �?        UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?      �?        �������?UUUUUU�?      �?      �?      �?              �?              �?        T�n�W�?ï�Dz��?'u_[�?�V'u�?��VC��?�H%�e�?______�?�?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ��N��N�?�؉�؉�?      �?        <<<<<<�?�?ffffff�?333333�?      �?      �?      �?      �?      �?              �?      �?              �?      �?        �]�ڕ��?��+Q��?��[��[�?�A�A�?�Kh/��?h/�����?O��N���?;�;��?]t�E�?F]t�E�?      �?      �?      �?              �?                      �?      �?              �?      �?              �?      �?        O�;���?�RKE,�?SJ)��R�?��Zk���?              �?\��[���?�i�i�?8��18�?������?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?      �?      �?              �?        ������?Cy�5��?pX���o�?A��)A�?���,d!�?8��Moz�?      �?        �������?UUUUUU�?�$I�$I�?۶m۶m�?�m۶m��?�$I�$I�?۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?�$I�$I�?�m۶m��?              �?      �?      �?��y��y�?�a�a�?      �?        �?�?      �?        �������?�������?      �?      �?      �?              �?              �?      �?              �?;�;��?;�;��?vb'vb'�?;�;��?      �?                      �?      �?              �?      �?�������?�������?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ%�[6hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       R                    �?��l�Qf�?�           8�@                                    @0`�#��?�             n@                                  @�d���Ҹ?U             a@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?5�wAd�?S            �`@                                0Cd=@���.�6�?             G@        	       
                 03[:@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     C@                                   �?`���i��?5             V@                                 �=@@9G��?            �H@                                 �9@ 	��p�?             =@        ������������������������       �                     @                                   �?�C��2(�?             6@       ������������������������       �                     2@                                  �?@      �?             @        ������������������������       �                     �?                                   D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                    �C@               I                 `f7@      �?A             Z@              D                  �2@�{��?3            �T@                                  @X3_��?.            �Q@        ������������������������       �                     @               A                    �?      �?+             P@              0                    �?�m����?(            �M@               '                    �?���Q��?             D@       !       &                    �?�<ݚ�?             2@       "       #                 �|�9@      �?             0@        ������������������������       �                      @        $       %                 ���@؇���X�?
             ,@        ������������������������       �                      @        ������������������������       �        	             (@        ������������������������       �                      @        (       /                 ��&@�eP*L��?             6@       )       .                    �?�q�q�?
             2@       *       +                 ���@      �?	             0@        ������������������������       �                     @        ,       -                    3@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     @        1       @                    �?�����?             3@       2       ?                    @ҳ�wY;�?             1@       3       4                 �!@     ��?             0@        ������������������������       �                     �?        5       6                   �,@������?             .@        ������������������������       �                     �?        7       :                    �?d}h���?
             ,@        8       9                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ;       <                 �|�;@�����H�?             "@       ������������������������       �                     @        =       >                 �|Y>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        B       C                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        E       F                 ���4@�C��2(�?             &@       ������������������������       �                     @        G       H                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        J       M                    @��2(&�?             6@        K       L                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        N       O                 ��T?@�}�+r��?             3@        ������������������������       �                     $@        P       Q                 ��p@@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        S       �                 ��D:@z�G�z�?.           `}@       T       �                    �?      �?�            �u@       U       �                    �?P9<h�;�?�            �s@       V       W                 ���@4��?�?�            �s@        ������������������������       �                     @@        X       Y                 ��@ �Cc}�?�            �q@        ������������������������       �                     �?        Z       o                   @4@����?�            pq@        [       \                     @V������?            �B@        ������������������������       �                     @        ]       ^                   �0@�!���?             A@        ������������������������       �                     �?        _       `                    �?:ɨ��?            �@@        ������������������������       �                      @        a       n                 ��Y @r֛w���?             ?@       b       c                   �2@�ՙ/�?             5@        ������������������������       �                     @        d       g                   �3@�E��ӭ�?             2@       e       f                 �?�@�q�q�?             (@       ������������������������       �                     @        ������������������������       �և���X�?             @        h       i                 P�@r�q��?             @        ������������������������       �                     @        j       m                 @3�@�q�q�?             @       k       l                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        p       �                     @\����?�            @n@        q       r                    �?      �?             H@        ������������������������       �                      @        s       t                 �|Y=@��(\���?             D@        ������������������������       �        
             (@        u       v                 �|�=@ �Cc}�?             <@        ������������������������       �                     �?        w       �                    F@�>����?             ;@       x       y                   �'@�KM�]�?             3@        ������������������������       �                     @        z       �                    �?؇���X�?             ,@       {       |                    @@r�q��?             (@        ������������������������       �                     @        }       ~                   @A@      �?              @        ������������������������       �                     �?               �                   �3@؇���X�?             @       �       �                   @D@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?lW3�kC�?z            @h@        �       �                 ��$1@��� ��?%             O@       �       �                 �� @�^����?#            �M@       �       �                 ���@L紂P�?            �I@        �       �                   �7@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                    �?r�q��?             B@        �       �                   �<@d}h���?	             ,@        ������������������������       �                     @        �       �                   @@�z�G��?             $@       ������������������������       ��q�q�?             @        �       �                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                  ��@��2(&�?             6@        ������������������������       �                     @        �       �                 �|Y=@@�0�!��?
             1@        ������������������������       �                     @        ������������������������       �        	             ,@        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��) @�5[|/��?U            �`@       �       �                 �?�@�x�E~�?:            @V@       ������������������������       �        $            �J@        �       �                 �|Y>@�X�<ݺ?             B@       ������������������������       �                     7@        �       �                   �?@8�Z$���?	             *@        ������������������������       �                     �?        �       �                 @3�@�8��8��?             (@        �       �                   �A@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    ?@X�EQ]N�?            �E@       �       �                    �?�חF�P�?             ?@       �       �                 pf� @�+$�jP�?             ;@        ������������������������       �                     �?        �       �                 �|�=@8�Z$���?             :@       �       �                    (@�8��8��?             8@       �       �                   �;@�r����?	             .@        �       �                    9@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���"@�C��2(�?             &@        ������������������������       �                     @        �       �                   �<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    )@�5��?             ;@        ������������������������       �                     $@        �       �                 `v�1@�IєX�?
             1@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        �                          @�D����?Q            �_@       �       	                   �?�;_��?F            @\@       �       �                    �?X�Emq�?B            �Z@        �       �                   �H@�eP*L��?            �@@       �       �                   �1@���Q��?             >@        ������������������������       �                     @        �       �                 p"�X@��
ц��?             :@       �       �                    �?�q�q�?             2@       �       �                   �A@��
ц��?	             *@       �       �                 �|Y<@�z�G��?             $@        ������������������������       �                     @        �       �                   @@@և���X�?             @       �       �                 �|�=@���Q��?             @       �       �                 ��2>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?              @       �       �                    �?�q�q�?             @        ������������������������       �                      @        �       �                    �?      �?             @       �       �                    >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 03k:@b1<+�C�?,            @R@        ������������������������       �                     @        �       �                   �A@X�Cc�?+            �Q@        �       �                 0�E@      �?             <@        ������������������������       �                      @        �       �                 `fFJ@��Q��?             4@        ������������������������       �                     @        �       �                    �?     ��?	             0@       �       �                    �?�q�q�?             @       �       �                 �|�>@���Q��?             @       �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 `f�N@ףp=
�?             $@        ������������������������       �                      @        �       �                 ��-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                        )?@�����?             E@        �                          �?d}h���?             ,@       �                         @=@      �?	             (@       �                       `f�;@"pc�
�?             &@       �                          �J@z�G�z�?             $@        �       �                    H@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                               x#J@h�����?             <@        ������������������������       �                     0@                              `�iJ@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        
                         �?����X�?             @                               �G@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������}<����?�/���?�
V�
V�?X}*X}*�?�uy)�?�h�?n]�?UUUUUU�?UUUUUU�?              �?      �?        �rv��?֘HT��?Y�B��?���7���?      �?      �?              �?      �?                      �?F]t�E�?F]t�E�?9/���?������?�{a���?������?              �?F]t�E�?]t�E�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?������?��18�?��V��?{2~�ԓ�?              �?      �?      �?�V'u�?��}ylE�?�������?333333�?�q�q�?9��8���?      �?      �?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?        t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?      �?              �?�؉�؉�?;�;��?              �?      �?                      �?              �?Q^Cy��?^Cy�5�?�������?�������?      �?      �?              �?wwwwww�?�?              �?I�$I�$�?۶m۶m�?333333�?�������?      �?                      �?�q�q�?�q�q�?      �?              �?      �?              �?      �?                      �?      �?        333333�?�������?      �?                      �?F]t�E�?]t�E�?              �?�������?�������?              �?      �?        ��.���?t�E]t�?UUUUUU�?UUUUUU�?      �?                      �?�5��P�?(�����?      �?        �q�q�?�q�q�?              �?      �?        �������?�������?      �?      �?����?-hk�׹?�N��N��?ى�؉��?      �?        %I�$I��?۶m۶m�?              �?�ru���?�ojT���?�g�`�|�?o0E>��?      �?        �������?�������?              �?N6�d�M�?e�M6�d�?              �?���{��?�B!��?�<��<��?�a�a�?              �?�q�q�?r�q��?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        ���|���?"pc�
�?      �?      �?      �?        �������?333333�?      �?        %I�$I��?۶m۶m�?              �?�Kh/��?h/�����?�k(���?(�����?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?              �?      �?              �?۶m۶m�?�$I�$I�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?        �fy���?��4l7˳?�{����?�B!��?u_[4�?W'u_�?�������?�������?�������?�?              �?      �?        �������?UUUUUU�?I�$I�$�?۶m۶m�?      �?        ffffff�?333333�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?        ��.���?t�E]t�?      �?        ZZZZZZ�?�������?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        N6�d�M�?'�l��&�?����G�?p�\��?      �?        ��8��8�?�q�q�?      �?        ;�;��?;�;��?              �?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?      �?      �?              �?        w�qG�?qG�wĽ?�Zk����?��RJ)��?/�����?B{	�%��?              �?;�;��?;�;��?UUUUUU�?UUUUUU�?�������?�?      �?      �?      �?                      �?]t�E�?F]t�E�?      �?        �������?�������?      �?                      �?      �?                      �?      �?              �?        333333�?�������?              �?      �?        h/�����?/�����?              �?�?�?      �?      �?              �?      �?              �?        �0�0�?z��y���?��Ź��?�(�u���?5�x+��?�}�	��?]t�E�?t�E]t�?�������?333333�?              �?�؉�؉�?�;�;�?UUUUUU�?UUUUUU�?�؉�؉�?�;�;�?333333�?ffffff�?              �?۶m۶m�?�$I�$I�?333333�?�������?      �?      �?              �?      �?              �?                      �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        �;w�ܹ�?Ĉ#F��?              �?%I�$I��?�m۶m��?      �?      �?              �?ffffff�?�������?      �?              �?      �?UUUUUU�?UUUUUU�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?�������?              �?      �?      �?              �?      �?        =��<���?�a�a�?I�$I�$�?۶m۶m�?      �?      �?/�袋.�?F]t�E�?�������?�������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�	3 hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM#hjh))��}�(h,h/h0M#��h2h3h4hph<�h=Kub������       �                 `fK@�3)0�F�?�           8�@              k                     @4�^��\�?v           x�@                                  �8@A�b��?�            �l@                                   �?�c�����?!            �J@                               �܅4@|��?���?             ;@                                 �1@ҳ�wY;�?             1@        ������������������������       �                     @                                   �?8�Z$���?
             *@        	       
                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   &@�C��2(�?             &@                                  �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@                                   �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     :@               j                    �?4��P8O�?k            �e@              ;                     �?�)m��{�?j            `e@               8                    �?*O���?.             R@              '                    �?:���W�?(            �M@                                �|�;@������?
             .@        ������������������������       �                     �?                                `f&;@d}h���?	             ,@        ������������������������       �                     �?               &                    �?8�Z$���?             *@              !                    �?"pc�
�?             &@                                    D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        "       #                   `=@؇���X�?             @        ������������������������       �                     @        $       %                 p�i@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        (       3                   �>@�zv�X�?             F@       )       *                    �?�5��?             ;@        ������������������������       �                     @        +       2                    R@r�q��?             8@       ,       -                 ��$:@      �?             6@        ������������������������       �                      @        .       1                 `fF<@d}h���?	             ,@       /       0                    J@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        4       7                   �B@�IєX�?
             1@        5       6                 �TaA@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        9       :                    �?�n_Y�K�?             *@        ������������������������       �                     @        ������������������������       �                      @        <       Q                   @4@r٣����?<            �X@       =       P                    �?V��z4�?$             O@       >       G                    �?�̚��?#            �N@        ?       @                   �B@���N8�?             5@       ������������������������       �        	             ,@        A       F                   �J@����X�?             @       B       C                   �'@      �?             @        ������������������������       �                     �?        D       E                   �*@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        H       I                    �?P���Q�?             D@        ������������������������       �                     @        J       O                 �|�=@�X�<ݺ?             B@        K       L                   �'@r�q��?             (@       ������������������������       �                     @        M       N                 �|Y<@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     8@        ������������������������       �                     �?        R       [                    �?$G$n��?            �B@        S       X                    �?"pc�
�?             &@       T       W                   �B@؇���X�?             @        U       V                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        Y       Z                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        \       e                    �?ȵHPS!�?             :@       ]       d                    :@���}<S�?             7@       ^       c                   �C@r�q��?             (@       _       b                    �?�C��2(�?             &@        `       a                    <@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        f       g                    =@�q�q�?             @        ������������������������       �                     �?        h       i                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        l       �                    �? ��@��?�            �v@       m       �                    �?�uw\l��?�            pq@        n       u                    �?P�t��?0            @R@        o       t                    �?���N8�?             5@        p       q                 �|�5@      �?             @        ������������������������       �                      @        r       s                 ��%@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        v       �                    �?D>�Q�?             J@       w       �                 �|Y=@d}h���?             <@        x                           �?�q�q�?             "@       y       ~                   �9@      �?              @       z       {                 ���@���Q��?             @        ������������������������       �                     �?        |       }                   �5@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     3@        �       �                   `3@      �?             8@       �       �                 �|Y=@�C��2(�?             6@        �       �                  ��@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 03�@�X�<ݺ?	             2@        ������������������������       �                      @        �       �                   @'@      �?             0@       ������������������������       ���S�ۿ?             .@        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    %@LX�
]�?�            �i@        ������������������������       �                     �?        �       �                    �?�p ��?�            �i@        �       �                   �4@�g�y��?             ?@        �       �                   �3@�z�G��?             $@       �       �                 `F�+@և���X�?             @       �       �                   �2@      �?             @       �       �                 P��@�q�q�?             @        ������������������������       �                     �?        �       �                 ��!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @B@�ՙ/�?             5@       �       �                   P&@�����?             3@       �       �                    �?և���X�?
             ,@       �       �                  S�"@�n_Y�K�?	             *@       �       �                 ��� @�q�q�?             (@       �       �                    8@���Q��?             $@        ������������������������       �                     @        �       �                 �&B@z�G�z�?             @        ������������������������       �                     @        �       �                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?����?n            �e@       �       �                 �?�@ĴF���?g            �d@        �       �                 �|Y=@xL��N�?3            �R@       ������������������������       �                    �D@        �       �                 ��@�C��2(�?            �@@        ������������������������       �                     ,@        �       �                   �@�S����?             3@        �       �                 �|Y>@���Q��?             @        ������������������������       �                      @        �       �                 �&B@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                 @3�@,sI�v�?4            �V@        �       �                    :@      �?              @        ������������������������       �                     @        �       �                   �?@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 `�X#@������?0            �T@       �       �                   �0@��� ��?'             O@        ������������������������       �      �?             @        �       �                   �:@4և����?%             L@        ������������������������       �                     5@        �       �                    <@؇���X�?            �A@        ������������������������       �                     �?        �       �                 ���"@�t����?             A@       �       �                 ��) @(;L]n�?             >@       ������������������������       �                     3@        �       �                 ��y @�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             4@        ������������������������       �                     $@        �       �                    �?<�\`*��?4             U@       �       �                 �A7@X�<ݚ�?            �F@       �       �                    �?և���X�?            �A@        �       �                    �?�θ�?	             *@       �       �                    �?      �?             (@        �       �                    &@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���.@      �?              @       �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 P��%@�eP*L��?             6@        ������������������������       �                     @        �       �                    @@X�<ݚ�?             2@       �       �                    (@r�q��?             (@       ������������������������       �                     @        �       �                   �=@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?�θ�?            �C@        �       �                    @      �?             @       �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �̼6@b�h�d.�?            �A@        �       �                   �1@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?@4և���?             <@       �       �                 ��T?@�8��8��?             8@       ������������������������       �                     3@        �       �                 ��p@@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       "                   @      �?E             ^@       �       �                    �?��mo*�?C            �]@       ������������������������       �        %            �P@               !                   @��
ц��?             J@                                 �?      �?             H@                                �?��
ц��?            �C@                                �?X�<ݚ�?             ;@                             �̾w@��.k���?	             1@             
                �|Y<@�q�q�?             (@             	                  �9@      �?              @                               �4@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                              p"�X@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @                                 �?      �?	             (@                                �?�eP*L��?             &@                               �D@X�<ݚ�?             "@                                �?�q�q�?             @                                >@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                  @�q�q�?             "@        ������������������������       �                     @                              �|�;@���Q��?             @        ������������������������       �                      @                               �|�>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0M#KK��h2h3h4hVh<�h=Kub������������Rl���?�[�'��?e
�d�?5���7��?�,�����?-����b�?:�&oe�?�V�9�&�?	�%����?{	�%���?�������?�������?              �?;�;��?;�;��?      �?      �?              �?      �?        ]t�E�?F]t�E�?      �?      �?              �?      �?              �?        �������?�������?              �?      �?                      �?iȹ�. �?-o�`���?Kj+����?j+�����?�q�q�?�q�q�?_[4��?A�Iݗ��?wwwwww�?�?              �?I�$I�$�?۶m۶m�?              �?;�;��?;�;��?/�袋.�?F]t�E�?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?        ��.���?�袋.��?/�����?h/�����?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        ۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�?�?۶m۶m�?�$I�$I�?      �?                      �?      �?        ;�;��?ى�؉��?              �?      �?        >���>�?|���?2�c�1�?�s�9��??�%C���?�u�y���?��y��y�?�a�a�?              �?�m۶m��?�$I�$I�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ffffff�?�������?      �?        ��8��8�?�q�q�?�������?UUUUUU�?      �?        333333�?�������?      �?                      �?      �?                      �?к����?���L�?/�袋.�?F]t�E�?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?              �?      �?              �?      �?        ��N��N�?�؉�؉�?ӛ���7�?d!Y�B�?�������?UUUUUU�?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?mo�<~'�?KBfb�?y�G�?�n���?�4iҤI�?˖-[�l�?�a�a�?��y��y�?      �?      �?              �?      �?      �?              �?      �?                      �?b'vb'v�?vb'vb'�?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?333333�?�������?      �?              �?      �?              �?      �?                      �?              �?      �?              �?      �?]t�E�?F]t�E�?      �?      �?      �?                      �?��8��8�?�q�q�?      �?              �?      �?�������?�?      �?              �?      �?      �?                      �?�@*9/�?���VC�?              �?Q��+Q�?��+Q��?��{���?�B!��?ffffff�?333333�?�$I�$I�?۶m۶m�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?              �?        �a�a�?�<��<��?^Cy�5�?Q^Cy��?۶m۶m�?�$I�$I�?ى�؉��?;�;��?UUUUUU�?UUUUUU�?�������?333333�?              �?�������?�������?      �?              �?      �?              �?      �?                      �?      �?              �?                      �?      �?        ��֡�l�?/�I���?E�JԮD�?ە�]�ڵ?>�S��?L�Ϻ��?      �?        ]t�E�?F]t�E�?      �?        (������?^Cy�5�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        l�l��?��I��I�?      �?      �?      �?        �������?333333�?              �?      �?        �|����?������?�{����?�B!��?      �?      �?I�$I�$�?�m۶m۶?      �?        ۶m۶m�?�$I�$I�?              �?<<<<<<�?�?�������?�?      �?        ]t�E�?F]t�E�?              �?      �?              �?      �?              �?      �?              �?              �?        =��<���?�a�a�?r�q��?�q�q�?۶m۶m�?�$I�$I�?�؉�؉�?ى�؉��?      �?      �?      �?      �?              �?      �?              �?      �?      �?      �?      �?                      �?              �?              �?t�E]t�?]t�E�?      �?        �q�q�?r�q��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ى�؉��?�؉�؉�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?;��:���?_�_��?۶m۶m�?�$I�$I�?              �?      �?        n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        333333�?�������?              �?      �?              �?              �?      �?W'u_�?�<�"h�?              �?�;�;�?�؉�؉�?      �?      �?�؉�؉�?�;�;�?�q�q�?r�q��?�?�������?UUUUUU�?UUUUUU�?      �?      �?�������?�������?              �?      �?                      �?      �?                      �?�������?333333�?              �?      �?              �?      �?]t�E�?t�E]t�?r�q��?�q�q�?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������                           @�_%����?�           8�@               	                    @�3Ea�$�?             G@                                   �?�X�<ݺ?             B@                                   �?����X�?             @        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     =@        
                           @�z�G��?             $@        ������������������������       �                     @                                   @և���X�?             @        ������������������������       �                     �?                                   @      �?             @                                  �?      �?             @        ������������������������       �                      @                                ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @               �                  x#J@�[�^��?�           Ȅ@              _                  �#@�J�j�?d           H�@               *                    �?��ti�?�            @l@               !                 �|Y;@P����?             C@                               �?@�\��N��?             3@        ������������������������       �                     @                                    @�	j*D�?             *@                                  �?"pc�
�?
             &@                                  �?ףp=
�?	             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        "       '                    �?���y4F�?             3@       #       $                 ���@��S�ۿ?
             .@        ������������������������       �                     @        %       &                    �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        (       )                 ��� @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        +       @                   �8@�*/�8V�?�            �g@        ,       1                    �?z�G�z�?&             I@        -       .                 ��y@���Q��?             @        ������������������������       �                     �?        /       0                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        2       9                 �?�@���V��?#            �F@       3       8                 ���@ �q�q�?             8@        4       5                    6@      �?             @        ������������������������       �                     �?        6       7                 �&b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@        :       ?                    �?����X�?             5@       ;       >                 ��Y @r�q��?             2@        <       =                   �2@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             (@        ������������������������       �                     @        A       ^                    �?D��*�4�?[            @a@       B       K                    �?`�bV��?X            �`@        C       H                 03s@�X�<ݺ?             B@       D       E                  ��@      �?             @@       ������������������������       �                     4@        F       G                 �|Y=@�8��8��?	             (@        ������������������������       �                     �?        ������������������������       �                     &@        I       J                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        L       W                   �?@DE�SA_�??            @X@       M       R                 �|�=@�y��*�?&             M@       N       O                 ��) @ �h�7W�?#            �J@       ������������������������       �                    �E@        P       Q                 pf� @�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        S       V                 �̌!@z�G�z�?             @       T       U                   �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        X       Y                   @C@ ���J��?            �C@       ������������������������       �                     6@        Z       [                      @�IєX�?             1@        ������������������������       �                      @        \       ]                    D@��S�ۿ?
             .@        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                     @        `       �                 03#?@Х��L�?�            pt@       a       z                     �?~#M����?�            `p@        b       o                   �F@#z�i��?            �D@        c       d                    <@�㙢�c�?             7@        ������������������������       �                     @        e       f                    �?      �?             0@        ������������������������       �                     @        g       h                 �|Y=@�q�q�?             (@        ������������������������       �                     �?        i       n                    �?���!pc�?             &@       j       k                  Y>@z�G�z�?             $@       ������������������������       �                     @        l       m                  �>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        p       q                    �?X�<ݚ�?             2@        ������������������������       �                     �?        r       s                    �?��.k���?
             1@        ������������������������       �                     @        t       y                    R@X�Cc�?             ,@       u       x                    K@      �?             (@       v       w                   �G@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        {       �                    �?�:тr��?�            �k@        |       �                     @
;&����?             G@        }       �                    �?������?
             .@        ~                           �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�P�*�?             ?@        �       �                    �?������?             .@       �       �                    �?�q�q�?             (@        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @     ��?             0@       �       �                    @X�Cc�?	             ,@       �       �                    �?�	j*D�?             *@       ������������������������       �                      @        �       �                   `3@z�G�z�?             @        ������������������������       �                     @        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?B0�8���?l            �e@        �       �                    @���Q��?1             T@       �       �                    '@�n_Y�K�?0            �S@        �       �                    �?r�q��?             @        �       �                    "@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?ޚ)�?,             R@       �       �                 м�9@���e��?(            �P@       �       �                 �|Y=@~|z����?            �J@        �       �                 `f�)@�q�q�?             8@        �       �                    �?�z�G��?             $@       ������������������������       �                     @        �       �                   �&@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    /@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        �       �                     @8^s]e�?             =@       �       �                   �*@      �?
             0@       �       �                   �'@����X�?             ,@        �       �                   �J@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �A@      �?              @       ������������������������       �                     @        �       �                    D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�n_Y�K�?             *@        ������������������������       �                      @        �       �                     @�eP*L��?             &@       �       �                 ���.@X�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?����X�?             @       �       �                 ��1@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     @        ������������������������       �                      @        �       �                    #@��s��?;            �W@        ������������������������       �                      @        �       �                    �?����D��?9            @W@       �       �                    &@��ɉ�?%            @P@        �       �                     @�8��8��?	             (@       �       �                    5@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        �       �                   �*@�O4R���?            �J@       �       �                 �|�=@�g�y��?             ?@        �       �                   �(@$�q-�?	             *@        ������������������������       �                      @        �       �                 �|Y<@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �        	             2@        ������������������������       �        
             6@        ������������������������       �                     <@        �       �                    �?z�G�z�?(            @P@        �       �                    @      �?             6@       �       �                     @b�2�tk�?             2@       ������������������������       �                     $@        �       �                 ��p@@      �?              @        �       �                 ��T?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�<@ �#�Ѵ�?            �E@        �       �                     �?8�Z$���?             *@        �       �                 `f�D@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     >@        �                          @d}h���?H             \@       �       	                    �?�J��g��?E            �Z@       �       �                    �?�J�4�?@             Y@       ������������������������       �        ,            @Q@        �                         �H@�g�y��?             ?@       �       �                    �?�LQ�1	�?             7@        �       �                    �?�q�q�?             @       �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    6@ҳ�wY;�?
             1@        ������������������������       �                      @        �                          �?������?             .@       �                          @H@ףp=
�?             $@        ������������������������       �                     @                                 �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                 C@���Q��?             @                                >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        
                        �6@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������z���� �?@Bx��?��,d!�?����7��?�q�q�?��8��8�?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?              �?ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?      �?      �?              �?      �?      �?      �?                      �?      �?        J@����?l}����?^-n����?D�#{��?��|٠�?�ɗ�|�?Q^Cy��?�P^Cy�?�5��P�?y�5���?              �?vb'vb'�?;�;��?/�袋.�?F]t�E�?�������?�������?              �?      �?                      �?              �?(������?6��P^C�?�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?r1����?m�w6�;�?�������?�������?�������?333333�?      �?              �?      �?              �?      �?        [�[��?�>�>��?�������?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �m۶m��?�$I�$I�?�������?UUUUUU�?      �?      �?              �?      �?              �?                      �?ہ�v`��?)�3J���?��f��?�3�τ?�?��8��8�?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        ���_\�?����?�4�rO#�?GX�i��?��sHM0�?"5�x+��?      �?        ffffff�?333333�?              �?      �?        �������?�������?      �?      �?      �?                      �?              �?��-��-�?�A�A�?      �?        �?�?      �?        �������?�?              �?      �?              �?        `J�+���?AkQ���?DP{k�?w�_�	)�?ە�]���?�+Q��?d!Y�B�?�7��Mo�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        t�E]t�?F]t�E�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        r�q��?�q�q�?      �?        �������?�?              �?%I�$I��?�m۶m��?      �?      �?      �?      �?      �?                      �?      �?                      �?u��t���?QQ�?�Mozӛ�?Y�B��?�?wwwwww�?�������?�������?              �?      �?        �������?333333�?              �?      �?        �RJ)���?�Zk����?wwwwww�?�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?�m۶m��?%I�$I��?;�;��?vb'vb'�?              �?�������?�������?      �?              �?      �?              �?      �?              �?              �?        �JC�}�?��jyc�?�������?333333�?ى�؉��?;�;��?�������?UUUUUU�?      �?      �?              �?      �?              �?        ��8��8�?9��8���?>���>�?�>���?��sHM0�?�	�[���?UUUUUU�?UUUUUU�?333333�?ffffff�?              �?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?              �?      �?        	�=����?|a���?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?ى�؉��?;�;��?              �?]t�E�?t�E]t�?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?                      �?              �?      �?        q�����?�X�0Ҏ�?              �?P?���O�?X`��??�?��? �����?UUUUUU�?UUUUUU�?]t�E�?F]t�E�?              �?      �?              �?        :�&oe�?�x+�R�?��{���?�B!��?�؉�؉�?;�;��?      �?        ]t�E�?F]t�E�?      �?                      �?      �?              �?              �?        �������?�������?      �?      �?9��8���?�8��8��?              �?      �?      �?      �?      �?      �?                      �?      �?              �?        �/����?�}A_Ч?;�;��?;�;��?      �?      �?              �?      �?              �?              �?        ۶m۶m�?I�$I�$�?�#蝺�?7��XQ�?{�G�z�?�z�G��?              �?�B!��?��{���?d!Y�B�?Nozӛ��?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?        �������?�������?      �?        �?wwwwww�?�������?�������?              �?UUUUUU�?�������?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ۶m۶m�?�$I�$I�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��~hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                  x#J@�C��ӽ�?�           8�@                                  @�P�2�?i           P�@                                   �?z�G�z�?             D@                                  @$�q-�?             :@       ������������������������       �                     8@        ������������������������       �                      @                                   �?X�Cc�?             ,@        ������������������������       �                     @        	                           �?      �?             $@        
                           @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   @      �?              @                                  @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               S                 ���"@rA3��k�?S           �@               "                    �?�jt����?�            �m@                                   �?�z�G��?             D@       ������������������������       �                     8@               !                 �|Y>@      �?
             0@                               pf�@z�G�z�?	             .@                                �|Y:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  �9@�8��8��?             (@       ������������������������       �                     @                                �?�@z�G�z�?             @        ������������������������       �                      @                                 @3�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        #       ,                    �?��A9G�?            �h@        $       +                 �|Y=@������?             A@        %       *                   �<@և���X�?             ,@       &       )                   �6@      �?              @        '       (                 ��y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     4@        -       2                    �?�X�<ݺ?j            @d@        .       /                  ��@�nkK�?             7@        ������������������������       �                     @        0       1                 �|Y=@      �?
             0@        ������������������������       �                     �?        ������������������������       �        	             .@        3       R                    �?P����Ż?[            `a@       4       M                    �?�IєX�?Z             a@       5       6                     @ �#�Ѵ�?U             `@        ������������������������       �                     *@        7       D                 �|Y>@�8���?M             ]@       8       9                   �7@�d���?9            �U@        ������������������������       �                     C@        :       ?                   @8@@9G��?"            �H@        ;       >                 `fF@؇���X�?             @        <       =                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        @       C                 �?$@�Ń��̧?             E@        A       B                 ���@�8��8��?             (@       ������������������������       �                     @        ������������������������       �z�G�z�?             @        ������������������������       �                     >@        E       L                   @@@\-��p�?             =@        F       I                   �?@      �?              @        G       H                 pff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        J       K                 P�@      �?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        ������������������������       �                     5@        N       O                 P�@����X�?             @       ������������������������       �                     @        P       Q                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        T       �                    �?�������?�            `s@        U       p                     @�����?S            �`@       V       e                    �?��S�ۿ?,            �R@       W       b                    L@ �h�7W�?!            �J@       X       _                   �H@`'�J�?            �I@       Y       ^                 ��*@`���i��?             F@        Z       ]                   �9@ �q�q�?             8@        [       \                    5@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             1@        ������������������������       �                     4@        `       a                     �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        c       d                   �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        f       g                    �?�C��2(�?             6@        ������������������������       �                     @        h       i                     �?�r����?             .@        ������������������������       �                     �?        j       o                    �?؇���X�?             ,@       k       l                   �8@r�q��?             (@        ������������������������       �                     @        m       n                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        q       ~                 �|Y=@o����?'             M@       r       y                    �?     ��?             @@        s       v                    �?�q�q�?             @        t       u                    5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        w       x                    '@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        z       }                  �M$@ ��WV�?             :@        {       |                   �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@               �                 ��p@@�n_Y�K�?             :@       �       �                   �D@���N8�?             5@       �       �                    �?z�G�z�?             4@        �       �                 P�h2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?r�q��?             2@        ������������������������       �                     @        �       �                   �B@d}h���?	             ,@       �       �                   @B@      �?             (@       �       �                    �?"pc�
�?             &@       �       �                 03�1@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|Y>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    $@L(ݧa��?i             f@        �       �                   �<@      �?             (@        ������������������������       �                     @        �       �                   �?@�q�q�?             "@       �       �                 �|�=@؇���X�?             @       �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     �?�Uk���?c            �d@        �       �                    �?�3Ea�$�?             G@        �       �                 ��2>@�S����?	             3@        �       �                 �|�=@�q�q�?             "@        �       �                 �ܵ<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    R@�<ݚ�?             ;@       �       �                    �?      �?             8@       �       �                 `f�;@��2(&�?             6@        �       �                   �K@����X�?             @       �       �                 X�,@@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �<@��S�ۿ?
             .@        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                      @        ������������������������       �                     @        �       �                     @T(y2��?I            �]@       �       �                    �? ��PUp�?+            �Q@       �       �                 `f�)@����?�?            �F@        ������������������������       �                     *@        �       �                 �|�=@      �?             @@        �       �                 �|�<@@4և���?	             ,@       ������������������������       �                     (@        �       �                 ��,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     :@        �       �                 ��Y)@8��8���?             H@        ������������������������       �                      @        �       �                 �|�?@�q��/��?             G@       �       �                    9@�חF�P�?             ?@       �       �                    �?�X�<ݺ?             2@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                 ��-@�	j*D�?	             *@        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@       �       �                 �|�;@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   `3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             .@        �       �                    �?2]��a�?P            @_@       �       �                 ���Q@�nkK�?,            @Q@        �       �                 �|�=@�����H�?             2@       �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?���J��?!            �I@       ������������������������       �                    �F@        �       �                    '@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       
                   @~h����?$             L@       �                           �?D7�J��?#            �K@       �                          �?�eP*L��?             F@       �       �                    �?      �?             D@        �       �                   �8@��Q��?             4@        �       �                    �?����X�?             @        ������������������������       �                     @        �       �                 �nc@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    I@8�Z$���?	             *@       �       �                 X�,@@�8��8��?             (@        �       �                 Ȫ�c@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��Q��?             4@        ������������������������       �                     �?        �       �                 03�M@p�ݯ��?             3@        �       �                 `�iJ@և���X�?             @        ������������������������       �                     �?        �       �                 `f�K@      �?             @       �       �                    7@���Q��?             @        ������������������������       �                      @        �       �                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �                          �?      �?             (@       �                           �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @              	                �|�>@���!pc�?             &@                             p�O@�����H�?             "@                              �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub���������������sI,�?��m��?슍���?(���"��?ffffff�?ffffff�?;�;��?�؉�؉�?              �?      �?        �m۶m��?%I�$I��?              �?      �?      �?      �?      �?      �?                      �?      �?      �?�������?�������?              �?      �?              �?        �j��j��?3*�2*��?E�pR���?�<�"h�?333333�?ffffff�?              �?      �?      �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?N��)x9�?����>4�?xxxxxx�?�?۶m۶m�?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        ��8��8�?�q�q�?�Mozӛ�?d!Y�B�?      �?              �?      �?              �?      �?        =}���(�?4,�T�w�?�?�?�/����?�}A_Ч?      �?        j��FX�?a���{�?�:���C�?Ȥx�L��?      �?        ������?9/���?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        ��<��<�?�a�a�?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?        a����?�{a���?      �?      �?      �?      �?      �?                      �?      �?      �?              �?333333�?�������?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ;T�Cu;�?�W�x��?^Cy�5�?Q^Cy��?�?�������?"5�x+��?��sHM0�?�?�������?F]t�E�?F]t�E�?UUUUUU�?�������?�$I�$I�?۶m۶m�?              �?      �?                      �?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?      �?                      �?F]t�E�?]t�E�?              �?�?�������?              �?�$I�$I�?۶m۶m�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�FX�i�?5�rO#,�?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?      �?                      �?O��N���?;�;��?      �?      �?              �?      �?              �?        ى�؉��?;�;��?��y��y�?�a�a�?�������?�������?      �?      �?      �?                      �?UUUUUU�?�������?              �?۶m۶m�?I�$I�$�?      �?      �?F]t�E�?/�袋.�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?              �?        �C!����?�z���?      �?      �?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?        ��?����?`�1`�?����7��?��,d!�?(������?^Cy�5�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        9��8���?�q�q�?      �?      �?��.���?t�E]t�?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        �������?�?              �?      �?              �?                      �?�F��F��?�5�5�?��ۥ���?��V،?��I��I�?l�l��?      �?              �?      �?n۶m۶�?�$I�$I�?      �?              �?      �?              �?      �?              �?              �?        UUUUUU�?�������?              �?�B����?��Mozӻ?�Zk����?��RJ)��?��8��8�?�q�q�?      �?      �?      �?                      �?      �?        vb'vb'�?;�;��?      �?        r�q��?�q�q�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        ����Mb�?+����?d!Y�B�?�Mozӛ�?�q�q�?�q�q�?      �?      �?              �?      �?                      �?�?______�?              �?UUUUUU�?�������?      �?                      �?%I�$I��?�m۶m��?J��yJ�?k߰�k�?]t�E�?t�E]t�?      �?      �?ffffff�?�������?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?      �?                      �?      �?        �������?ffffff�?      �?        ^Cy�5�?Cy�5��?۶m۶m�?�$I�$I�?              �?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?                      �?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?      �?              �?      �?              �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM%hjh))��}�(h,h/h0M%��h2h3h4hph<�h=Kub������                         �R@>AU`�z�?�           8�@                                  @$5;Uʹ�?�            �@                                   @���N8�?             E@       ������������������������       �                     =@                                   @�θ�?	             *@        ������������������������       �                     @                                   �?      �?             @              	                    @      �?             @        ������������������������       �                     �?        
                           @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               c                    �?pTV�h�?�           Ђ@               6                 �|Y=@�Gi����?a            �b@                                 ��@��Q:��?#            �M@                                   �?�q�q�?             (@                                  �?X�<ݚ�?             "@        ������������������������       �                     �?                                   �?      �?              @                                 @9@և���X�?             @                               ��y@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                  P,@p�v>��?            �G@        ������������������������       �        	             3@                3                    �?      �?             <@       !       "                     �?�q�����?             9@        ������������������������       �                     @        #       ,                   �8@�����?             3@       $       %                    )@r�q��?             (@        ������������������������       �                     @        &       )                     @����X�?             @        '       (                 ��6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        *       +                    3@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        -       .                    �?և���X�?             @        ������������������������       �                     �?        /       0                     @      �?             @        ������������������������       �                      @        1       2                 �0@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        4       5                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        7       b                   �K@�ZD����?>            @V@       8       a                   @J@�J�j�?7            �S@       9       T                    �?���!pc�?6            @S@       :       M                    �?&����?,            @P@        ;       F                 ���4@؇���X�?            �A@       <       E                 X�@@`2U0*��?             9@       =       >                     @�}�+r��?             3@        ������������������������       �                      @        ?       D                    �?�IєX�?
             1@       @       C                   @@$�q-�?	             *@       A       B                 ���@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        G       L                   �F@���Q��?             $@       H       K                 �|�=@և���X�?             @        I       J                 ��2>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        N       S                    �?�z�G��?             >@        O       R                    �?      �?             (@       P       Q                  ��@ףp=
�?	             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     2@        U       V                     �?�q�q�?
             (@        ������������������������       �                      @        W       X                     @      �?	             $@        ������������������������       �                     �?        Y       `                    �?X�<ݚ�?             "@       Z       [                    �?և���X�?             @        ������������������������       �                      @        \       ]                    �?z�G�z�?             @        ������������������������       �                     �?        ^       _                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        d       �                    �?�� 27��?)           `|@        e       ~                     @�q�q�?V            �`@       f       }                    �?l��\��?.             Q@       g       v                  �v7@�p ��?            �D@        h       m                   �;@      �?             4@        i       l                    �?      �?             @       j       k                   �'@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        n       u                    L@      �?             0@       o       t                   �*@��S�ۿ?
             .@       p       q                   �'@�C��2(�?             &@        ������������������������       �                     �?        r       s                   �B@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        w       |                 `fF:@���N8�?             5@       x       y                    D@$�q-�?	             *@       ������������������������       �                      @        z       {                     �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ;@               �                 ���5@     ��?(             P@       �       �                    �?      �?             D@       �       �                    A@��>4և�?             <@       �       �                 ���@`�Q��?             9@        ������������������������       �                     @        �       �                 �|Y>@���|���?             6@       �       �                 �|Y<@D�n�3�?             3@       �       �                   �9@b�2�tk�?             2@       �       �                    �?     ��?	             0@       �       �                    7@��
ц��?             *@       �       �                    4@���Q��?             $@        �       �                 ��!@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �̜!@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�q�q�?             (@       �       �                 03�0@����X�?             @       �       �                 �|Y;@r�q��?             @        �       �                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �=@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �? �q�q�?             8@        �       �                    @�����H�?             "@        ������������������������       �                     @        �       �                   @C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        �       �                    �?Qv4@�?�             t@       �       �                 ��$:@�r����?�            �p@       �       �                   �0@�D�d@6�?�            �m@        �       �                 hf1@և���X�?             @       �       �                 pf�@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        �       �                   @A@�C��2(�?�            �l@       �       �                 �|�=@��CC`)�?t            �f@       �       �                 �|Y=@�J��_��?c            �c@       �       �                     @d����?E            �\@        �       �                    5@$�q-�?             :@        �       �                    &@r�q��?             (@        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �        
             ,@        �       �                   �<@xP�Fֺ�?5            @V@       �       �                   �:@�8��8��?3             U@       �       �                 ���@0z�(>��?-            �Q@        �       �                   �8@      �?              @       �       �                 ���@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@�i�y�?(            �O@       ������������������������       �                     C@        �       �                 0S5 @HP�s��?             9@        �       �                   �3@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     1@        �       �                   �;@�	j*D�?             *@        ������������������������       �                     @        ������������������������       �                     "@        �       �                 �̌!@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                  sW@`���i��?             F@        �       �                 pf�@�X�<ݺ?             2@       ������������������������       �        	             0@        ������������������������       �      �?              @        ������������������������       �                     :@        �       �                     @���!pc�?             6@        �       �                 `fF)@      �?              @       ������������������������       �                     @        �       �                    @@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �?@X�Cc�?
             ,@        �       �                   �>@      �?             @       �       �                 (Se!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �@z�G�z�?             $@        �       �                   �@@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �C@p���?             I@        �       �                 �?�@�IєX�?             1@        ������������������������       �                     @        �       �                   �B@ףp=
�?             $@        ������������������������       �                     �?        �       �                 ���$@�����H�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                    �@@        �       �                     �?      �?             @@       �       �                   �>@�5��?             ;@        �       �                    D@      �?	             (@        ������������������������       �                     @        �       �                   �Q@���Q��?             @       �       �                   @J@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|�<@�r����?	             .@        ������������������������       �                      @        ������������������������       �                     *@        �       �                     @z�G�z�?             @        ������������������������       �                     �?        �       �                    ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �                       ��9L@0G���ջ?&             J@       �                       ��l#@ qP��B�?!            �E@                               P�@r�q��?             @       ������������������������       �                     @                                 �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �B@                                  �?�<ݚ�?             "@                                >@���Q��?             @        ������������������������       �                      @        	      
                   P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?t�U����?-            �P@                              "�b@`Ql�R�?            �G@       ������������������������       �                     >@                                 !@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �        
             0@                                 �?��Q��?             4@                              �6f@���!pc�?             &@                               �5@z�G�z�?             $@        ������������������������       �                     �?                                �D@�����H�?             "@        ������������������������       �                     @                                 �?z�G�z�?             @        ������������������������       �                      @                              ���[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?              $                   �?X�<ݚ�?             "@              #                �̾w@և���X�?             @       !      "                `��`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0M%KK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?��6�?��2����?��y��y�?�a�a�?              �?ى�؉��?�؉�؉�?      �?              �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        ��O�?�̫�a��?o0E>��?#�u�)��?�A�I��?'u_[�?UUUUUU�?UUUUUU�?r�q��?�q�q�?              �?      �?      �?�$I�$I�?۶m۶m�?�������?333333�?      �?                      �?      �?              �?              �?        L� &W�?ڨ�l�w�?              �?      �?      �?�p=
ף�?���Q��?              �?Q^Cy��?^Cy�5�?�������?UUUUUU�?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        |��^���?	E(B��?^-n����?D�#{��?F]t�E�?t�E]t�?�����?�����?۶m۶m�?�$I�$I�?���Q��?{�G�z�?�5��P�?(�����?      �?        �?�?�؉�؉�?;�;��?۶m۶m�?�$I�$I�?      �?              �?      �?      �?              �?              �?        333333�?�������?۶m۶m�?�$I�$I�?      �?      �?              �?      �?                      �?      �?        ffffff�?333333�?      �?      �?�������?�������?      �?                      �?      �?              �?        �������?�������?              �?      �?      �?      �?        �q�q�?r�q��?�$I�$I�?۶m۶m�?              �?�������?�������?      �?              �?      �?      �?                      �?              �?              �?      �?        U���g�?W�N~0��?UUUUUU�?UUUUUU�?�������?------�?��+Q��?Q��+Q�?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?�?�������?F]t�E�?]t�E�?              �?�������?�������?              �?      �?                      �?      �?        �a�a�?��y��y�?;�;��?�؉�؉�?              �?�������?�������?              �?      �?                      �?              �?      �?      �?      �?      �?I�$I�$�?۶m۶m�?{�G�z�?��(\���?              �?F]t�E�?]t�E]�?(������?l(�����?9��8���?�8��8��?      �?      �?�;�;�?�؉�؉�?�������?333333�?      �?      �?      �?                      �?      �?      �?              �?      �?              �?                      �?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?�$I�$I�?�m۶m��?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?        �������?333333�?      �?                      �?�������?UUUUUU�?�q�q�?�q�q�?      �?              �?      �?              �?      �?              �?        �6��?̀O��?�������?�?}��|���?���й?�$I�$I�?۶m۶m�?�������?333333�?      �?              �?      �?      �?        ]t�E�?F]t�E�?�J�v�?4O��I�?d�^�.�?�%w��?�����a�?�(�j�?�؉�؉�?;�;��?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        �.p��?�я~���?UUUUUU�?UUUUUU�?�ԓ�ۥ�?H���@��?      �?      �?      �?      �?      �?                      �?      �?        �������?AA�?      �?        q=
ףp�?{�G�z�?      �?      �?              �?      �?              �?        vb'vb'�?;�;��?              �?      �?        �������?�������?      �?                      �?F]t�E�?F]t�E�?��8��8�?�q�q�?      �?              �?      �?      �?        F]t�E�?t�E]t�?      �?      �?      �?              �?      �?      �?                      �?%I�$I��?�m۶m��?      �?      �?      �?      �?      �?                      �?              �?�������?�������?      �?      �?              �?      �?              �?        \���(\�?{�G�z�?�?�?      �?        �������?�������?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?              �?              �?      �?h/�����?/�����?      �?      �?              �?333333�?�������?      �?      �?      �?      �?      �?                      �?�������?�?              �?      �?        �������?�������?      �?              �?      �?              �?      �?        vb'vb'�?�؉�؉�?��}A�?�}A_З?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        9��8���?�q�q�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        g��1��?���-�?W�+�ɕ?}g���Q�?              �?�?�?      �?                      �?ffffff�?�������?t�E]t�?F]t�E�?�������?�������?      �?        �q�q�?�q�q�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?r�q��?�$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?              �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�DhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       F                    �?��ϙLq�?�           8�@                                   �?D������?{            `h@                                    @���(`�?3            �U@       ������������������������       �                     K@                                   �?r٣����?            �@@              	                 ���@ȵHPS!�?             :@                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        
                        ���,@���}<S�?             7@       ������������������������       �        	             ,@                                 S�-@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @                                `�@1@����X�?             @        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               /                     �?\�f<t�?H             [@               .                    �?�ʻ����?             A@              -                    �?     ��?             @@              $                 ��UO@`՟�G��?             ?@              #                    �?����X�?             ,@                                Y>@�θ�?             *@                                �|�;@�q�q�?             @        ������������������������       �                     �?                                X�,@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               "                 p�i@@ףp=
�?             $@                !                  �>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        %       (                   �8@j���� �?             1@        &       '                 ���Q@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        )       *                 p"�X@z�G�z�?             $@       ������������������������       �                     @        +       ,                 p�w@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        0       E                    �?������?/            �R@       1       <                   �6@(N:!���?,            �Q@        2       7                   �2@���|���?             &@        3       4                    �?���Q��?             @        ������������������������       �                      @        5       6                 ��}@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        8       ;                    5@r�q��?             @       9       :                 �{@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        =       D                 �|�=@P����?%            �M@       >       ?                 �|=@��<b�ƥ?             G@        ������������������������       �                      @        @       A                    �?P�Lt�<�?             C@       ������������������������       �                    �A@        B       C                 ��.@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �                     @        G       �                     @BV�(��?G            �@        H       �                    �?o�����?�             m@       I       �                 `��R@���Q��?i            @e@       J       K                    @.���ڨ�?b            �c@        ������������������������       �                     @        L       �                   �K@,���y4�?^             c@       M       n                     �?h�wl�I�?U            �`@        N       m                   @I@և���X�?            �H@       O       P                    �?F�����?            �F@        ������������������������       �                     @        Q       l                   �H@�z�G��?             D@       R       c                    �?4�B��?            �B@       S       b                   �G@     ��?             @@       T       a                   �F@>���Rp�?             =@       U       \                   @@@�q�q�?             5@       V       [                   �>@      �?
             0@        W       X                 �|�<@և���X�?             @        ������������������������       �                     �?        Y       Z                 `fF<@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ]       ^                 03k:@���Q��?             @        ������������������������       �                     �?        _       `                   �C@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        d       k                 03�M@���Q��?             @       e       j                 `f�K@      �?             @       f       g                    7@�q�q�?             @        ������������������������       �                     �?        h       i                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        o       �                   �:@�ģ�a@�?6            @U@       p       w                    �?�o;����?3            �S@        q       r                   �2@(;L]n�?             >@       ������������������������       �                     4@        s       v                   �7@ףp=
�?             $@        t       u                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        x       {                    &@�q��/��?            �H@        y       z                   �5@�q�q�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        |       �                    �?��(\���?             D@       }       �                   �*@�C��2(�?            �@@       ~                        `fF)@�����H�?             ;@        ������������������������       �                      @        �       �                   @D@H%u��?             9@       ������������������������       �        	             1@        �       �                    G@      �?              @        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `fF<@�X�<ݺ?	             2@       ������������������������       �                     "@        �       �                   �Q@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|�=@�C��2(�?             &@        �       �                 �|Y=@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?r֛w���?+             O@       �       �                    �?^������?            �A@       ������������������������       �                     4@        �       �                    *@z�G�z�?             .@        ������������������������       �                     @        ������������������������       �                     (@        �       �                    @PN��T'�?             ;@       �       �                     �?ȵHPS!�?             :@        �       �                    @�����H�?             "@        �       �                 �(\�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�t����?
             1@        ������������������������       �                     "@        �       �                    �?      �?              @       �       �                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `fF6@$�`��S�?�            �q@       �       �                  �#@T�r�;�?�            �m@       �       �                    �?L���#��?p             f@       �       �                 ���@|T(W�j�?j            �d@        ������������������������       �                     ,@        �       �                   �2@L:�f@�?_            �b@        �       �                 ��@�	j*D�?	             *@       �       �                    �?      �?              @        �       �                 P��@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �0@���Q��?             @        ������������������������       �                     �?        �       �                 ��Y @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���@���}<S�?V            @a@        ������������������������       �                     �?        �       �                 �Yu@�<_���?U             a@        �       �                 P�N@      �?             D@       �       �                    7@l��\��?             A@        �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     :@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �?�@�*v��?>            @X@        ������������������������       �                     <@        �       �                 @3�@���}<S�?-            @Q@        �       �                    :@�q�q�?             "@        ������������������������       �                     @        �       �                   �?@      �?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        �       �                   �3@P���Q�?'             N@        �       �                 0S5 @      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        �       �                 ���"@h�����?$             L@       �       �                    <@p���?             I@        �       �                   �:@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                     >@        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                 �|�=@      �?             @        ������������������������       �                      @        �       �                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���!pc�?             &@       �       �                 P�@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    )@�ɞ`s�?)            �N@        �       �                     @�	j*D�?
             *@       ������������������������       �                     "@        ������������������������       �                     @        �       �                    �?�q�q�?             H@        �       �                    �?���Q��?             9@        �       �                    4@z�G�z�?             @        ������������������������       �                      @        �       �                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|Y=@�z�G��?             4@        ������������������������       �                     &@        �       �                   �D@�q�q�?             "@       �       �                     @؇���X�?             @       �       �                 03�1@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@        �       �                    �?`Ql�R�?            �G@        �       �                    @ ��WV�?             :@       ������������������������       �        
             4@        �       �                 ���A@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������Ӭ����?�X�>��?_�^��?�����?Ȥx�L��?g��o��?              �?|���?>���>�?�؉�؉�?��N��N�?UUUUUU�?UUUUUU�?              �?      �?        d!Y�B�?ӛ���7�?              �?�q�q�?9��8���?      �?                      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?��Kh/�?&���^B�?�������?<<<<<<�?      �?      �?�1�c��?�s�9��?�m۶m��?�$I�$I�?ى�؉��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?�������?�������?�������?      �?                      �?      �?                      �?ZZZZZZ�?�������?�m۶m��?�$I�$I�?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?              �?      �?        ��g�`��?к����?|�W|�W�?�A�A�?F]t�E�?]t�E]�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?�������?�������?      �?                      �?              �?�V'u�?'u_[�?��7��M�?d!Y�B�?      �?        ���k(�?(�����?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �/����?��/���?�i��F�?#,�4�r�?333333�?�������?g@(�S�?�1��X�?      �?        ������?����k�?T�n�Wc�?Xc"=P9�?�$I�$I�?۶m۶m�?�>�>��?؂-؂-�?              �?ffffff�?333333�?�Y7�"��?L�Ϻ��?      �?      �?�i��F�?GX�i���?UUUUUU�?UUUUUU�?      �?      �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?      �?        �������?333333�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?              �?                      �?rrrrrr�?�?�#{���?��	�Z�?�?�������?              �?�������?�������?      �?      �?              �?      �?                      �?/����?և���X�?UUUUUU�?UUUUUU�?      �?      �?      �?        �������?333333�?]t�E�?F]t�E�?�q�q�?�q�q�?      �?        )\���(�?���Q��?      �?              �?      �?�������?333333�?      �?              �?              �?        �������?UUUUUU�?              �?      �?        ��8��8�?�q�q�?      �?        �q�q�?�q�q�?      �?                      �?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?�B!��?���{��?_�_��?uPuP�?              �?�������?�������?              �?      �?        h/�����?&���^B�?�؉�؉�?��N��N�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?�?<<<<<<�?              �?      �?      �?�$I�$I�?�m۶m��?              �?      �?                      �?      �?        as �
��?{2~�ԓ�?��ǃ��?�Ӭ����?�.�袋�?��.�袻?��YΟ��?�0�Ӹ?      �?        �o�7���?ـl@6 �?vb'vb'�?;�;��?      �?      �?      �?      �?              �?      �?              �?        �������?333333�?              �?      �?      �?              �?      �?        ӛ���7�?d!Y�B�?              �?p�h�?n�?ܺ���?      �?      �?------�?�������?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        ���AG�? tT����?      �?        ӛ���7�?d!Y�B�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?333333�?�������?ffffff�?�������?      �?      �?      �?      �?      �?        �m۶m��?�$I�$I�?\���(\�?{�G�z�?ffffff�?�������?      �?                      �?      �?        �������?UUUUUU�?      �?              �?      �?      �?              �?      �?              �?      �?        F]t�E�?t�E]t�?      �?      �?              �?      �?              �?        mާ�d�?&C��6��?;�;��?vb'vb'�?              �?      �?        UUUUUU�?�������?333333�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?ffffff�?333333�?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?�������?              �?      �?                      �?      �?              �?        }g���Q�?W�+�ɕ?O��N���?;�;��?      �?        �������?UUUUUU�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���MhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       r                     @*�Ⱦ��?�           8�@               I                    �?�|@ߑ��?�            0t@              8                 ��UO@#F���?�            `k@              )                   �F@���Q��?j            �d@                                  �?p<�w���?N            �_@                                   �?$��m��?             :@                                  �?�\��N��?             3@        ������������������������       �                     @        	       
                 ���4@      �?	             (@        ������������������������       �                     @                                `f&;@�q�q�?             "@        ������������������������       �                     �?                                   �?      �?              @                               �|�;@����X�?             @        ������������������������       �                     �?                                   C@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?� �	��?>             Y@        ������������������������       �                    �A@               "                 `fF:@��ɉ�?)            @P@              !                   �D@�&=�w��?!            �J@                                   �? pƵHP�?              J@        ������������������������       �                     (@                                    �?�(\����?             D@                                 �@@ ���J��?            �C@       ������������������������       �                    �@@                                  @A@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        #       (                 X��B@�q�q�?             (@       $       '                   �<@      �?              @       %       &                 `f�D@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        *       /                 ���&@�ݜ�?            �C@        +       .                    �?���Q��?             @       ,       -                   �J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        0       1                 `fF:@l��\��?             A@        ������������������������       �        	             ,@        2       7                    K@R���Q�?             4@       3       6                 �T!@@�z�G��?             $@        4       5                   `G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        9       :                    �?�+$�jP�?             K@       ������������������������       �                     C@        ;       >                    �?      �?	             0@        <       =                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ?       @                 `��Q@�q�q�?             (@        ������������������������       �                      @        A       H                    �?z�G�z�?             $@       B       C                   �4@�q�q�?             @        ������������������������       �                     �?        D       G                    �?z�G�z�?             @       E       F                 �̾w@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        J       Y                    �?>�Q��?C             Z@       K       N                    @��S�ۿ?)             N@        L       M                     �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        O       T                   �E@���U�?'            �L@       P       S                    6@@��8��?              H@        Q       R                   �3@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     F@        U       V                    �?�����H�?             "@        ������������������������       �                     @        W       X                    G@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        Z       e                 `fFJ@�X���?             F@       [       \                    �?��2(&�?             6@       ������������������������       �                     ,@        ]       d                 �D C@      �?              @       ^       _                    �?����X�?             @        ������������������������       �                     @        `       a                   �2@      �?             @        ������������������������       �                     �?        b       c                    :@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        f       m                   �D@�eP*L��?             6@        g       h                    �?"pc�
�?             &@        ������������������������       �                     @        i       l                     �?      �?              @       j       k                    7@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        n       o                   �G@���!pc�?             &@        ������������������������       �                     @        p       q                   �L@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        s                          �?�j&|mH�?�            @x@       t                           /@��X��?�             u@        u       v                    #@���}<S�?             7@       ������������������������       �        
             (@        w       x                    &@"pc�
�?             &@        ������������������������       �                     �?        y       z                   �,@ףp=
�?             $@        ������������������������       �                     @        {       |                    �?z�G�z�?             @        ������������������������       �                      @        }       ~                   �-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�,�;i��?�            �s@        �       �                    �?*O���?.             R@        �       �                 X�,A@ �Cc}�?             <@       �       �                    �?�>����?             ;@       ������������������������       �                     5@        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �;@d�
��?             F@       �       �                    �?��H�}�?             9@       �       �                   �6@���y4F�?             3@       �       �                    3@�q�q�?             (@        �       �                   !@z�G�z�?             @        �       �                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                  p @և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 P�@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�d�����?             3@       �       �                 pf�$@�q�q�?             (@        ������������������������       �                     @        �       �                 03�1@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @@@:��A�?�             n@       �       �                    �?����f�?�            �h@        �       �                   �6@�f7�z�?             =@        �       �                 ��y@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             8@       �       �                    �?8����?             7@       �       �                 �|Y=@b�2�tk�?             2@        �       �                   �8@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���@�θ�?             *@        ������������������������       �                     @        �       �                 �|�=@�q�q�?             "@       �       �                   @@և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �>@��YIY�?o            �d@       �       �                 �|Y=@�v,D�?h            �c@       �       �                    �?��zi��?;            �V@        ������������������������       �                      @        �       �                    �?4\�����?:            @V@       �       �                 @3�@p#�����?3            �S@        ������������������������       �                     C@        �       �                   �<@���� �?            �D@       �       �                   �0@tk~X��?             B@        �       �                 �̌!@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                   �:@�חF�P�?             ?@       �       �                   �3@ȵHPS!�?             :@       �       �                   �1@     ��?	             0@        ������������������������       �                     @        �       �                   �2@�θ�?             *@        �       �                 ��Y @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 0S5 @�<ݚ�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �̌!@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�z�G��?             $@       �       �                 P�@      �?              @       ������������������������       �                     @        �       �                    6@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �Y5@t�e�í�?-            �P@        �       �                    �?�LQ�1	�?             7@       �       �                    �?��2(&�?             6@       �       �                 ���@��S�ۿ?             .@        ������������������������       �                     @        ������������������������       ������H�?             "@        �       �                 ��,@����X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     �?        �       �                 �|�=@���7�?             F@       �       �                    �?������?            �D@        ������������������������       �                     @        �       �                 ��) @ >�֕�?            �A@       ������������������������       �                     7@        �       �                 �̜!@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        �       �                 �&B@�q�q�?             "@        ������������������������       �                     �?        �       �                   �?@      �?              @        ������������������������       �                      @        �       �                 �!B@�q�q�?             @       �       �                 P�@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        �                          �?`Ӹ����?            �F@       �       �                    �?@-�_ .�?            �B@        ������������������������       �                     @        �       �                 �?�@`Jj��?             ?@        ������������������������       �        	             ,@        �       �                   @C@�t����?             1@        ������������������������       �                      @        �                         @D@�<ݚ�?             "@                               ��	0@�q�q�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                 @$�q-�?             J@             	                ���0@ףp=
�?             D@                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        
                         �?�IєX�?             A@                                 �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                 �?(;L]n�?             >@                              ��T?@��S�ۿ?             .@       ������������������������       �                     (@                              ��p@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                     (@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�����������������?�{d�_�?�X0��"�?��g?���?�������?+���?333333�?�������?!� ��?�������?vb'vb'�?�N��N��?�5��P�?y�5���?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?                      �?      �?                      �?�Q����?)\���(�?              �?�����?�����?tHM0���?�x+�R�?'vb'vb�?;�;��?      �?        333333�?�������?��-��-�?�A�A�?      �?        �������?UUUUUU�?              �?      �?              �?                      �?�������?�������?      �?      �?      �?      �?              �?      �?              �?                      �?\��[���?�i�i�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ------�?�������?      �?        333333�?333333�?ffffff�?333333�?      �?      �?      �?                      �?      �?              �?        B{	�%��?/�����?              �?      �?      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?      �?                      �?      �?              �?        ��N��N�?��؉���?�?�������?UUUUUU�?UUUUUU�?      �?                      �?p�}��?	�#����?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?�q�q�?�q�q�?              �?�������?�������?      �?                      �?]t�E�?�E]t��?��.���?t�E]t�?      �?              �?      �?�m۶m��?�$I�$I�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?]t�E�?t�E]t�?F]t�E�?/�袋.�?              �?      �?      �?�$I�$I�?۶m۶m�?      �?                      �?      �?        F]t�E�?t�E]t�?      �?        �������?333333�?              �?      �?        w�<�L��?���fy�?n۶m۶�?%I�$I��?d!Y�B�?ӛ���7�?              �?F]t�E�?/�袋.�?      �?        �������?�������?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?F܋��?u�G���?�q�q�?�q�q�?۶m۶m�?%I�$I��?h/�����?�Kh/��?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �袋.��?�.�袋�?
ףp=
�?{�G�z�?(������?6��P^C�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?                      �?�������?UUUUUU�?              �?      �?        Cy�5��?y�5���?�������?�������?      �?        UUUUUU�?�������?              �?      �?              �?        W�W��?��ƕ���?h�����?^N��)x�?O#,�4��?a���{�?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?d!Y�B�?8��Moz�?�8��8��?9��8���?�������?�������?      �?                      �?ى�؉��?�؉�؉�?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?�������?333333�?      �?              �?              �?                      �?��;���?��ұ�?~W��0��?�ґ=�?��_��_�?h�h��?              �?�{��^��?B�P�"�?7a~W��?�#{���?      �?        jW�v%j�?,Q��+�?r�q��?9��8���?333333�?�������?UUUUUU�?UUUUUU�?      �?        �Zk����?��RJ)��?��N��N�?�؉�؉�?      �?      �?      �?        ى�؉��?�؉�؉�?      �?      �?              �?      �?        9��8���?�q�q�?      �?      �?      �?              �?        333333�?�������?              �?      �?        �������?�������?      �?                      �?ffffff�?333333�?      �?      �?      �?              �?      �?              �?      �?              �?        �1����?�rv��?��Moz��?Y�B��?��.���?t�E]t�?�������?�?      �?        �q�q�?�q�q�?�m۶m��?�$I�$I�?      �?              �?      �?      �?        �.�袋�?F]t�E�?p>�cp�?������?      �?        ��+��+�?�A�A�?      �?        �������?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �??�>��?l�l��?S�n0E�?к����?      �?        ���{��?�B!��?      �?        <<<<<<�?�?      �?        9��8���?�q�q�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?              �?        �؉�؉�?;�;��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?        �?�?      �?      �?              �?      �?        �������?�?�������?�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ9M�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       Z                    �?\��m͗�?�           8�@                                03@r�=���?{            �h@                                   �?^l��[B�?#             M@                                ��y@�LQ�1	�?             7@        ������������������������       �                     �?                                   �?��2(&�?             6@        ������������������������       �                     �?               	                   @9@�����?             5@        ������������������������       �                     �?        
                        ���@P���Q�?             4@       ������������������������       �                     ,@                                �|=@r�q��?             @        ������������������������       �                      @        ������������������������       �      �?             @                                  �7@����X�?            �A@        ������������������������       �                     @                                �Y�@�n`���?             ?@                                   �?���|���?             &@                                ���@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   �?ףp=
�?             4@                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             0@               /                    �?Hg�m���?X            `a@              .                 03�=@ ����?-            @P@              -                    �?�'�`d�?            �@@              (                 �|Y=@p�ݯ��?             3@               !                    �?8�Z$���?
             *@        ������������������������       �                      @        "       '                 `�@1@���Q��?             @       #       $                    '@�q�q�?             @        ������������������������       �                     �?        %       &                   �,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        )       *                  S�2@r�q��?             @        ������������������������       �                     @        +       ,                      @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                     @@        0       Y                   �H@~�hP��?+            �R@       1       V                    C@p�EG/��?&            �O@       2       M                    �?���dQ'�?"            �L@       3       <                 ��5@p�v>��?            �G@        4       ;                    �?R���Q�?             4@       5       6                     @     ��?	             0@        ������������������������       �                     �?        7       :                 �|Y=@z�G�z�?             .@       8       9                 �&�)@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        =       L                    �?�5��?             ;@       >       ?                   �8@��H�}�?             9@        ������������������������       �                     @        @       A                    <@�G�z��?             4@        ������������������������       �                     @        B       E                 ��";@������?	             .@        C       D                     �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        F       G                 �|Y=@�C��2(�?             &@        ������������������������       �                      @        H       K                 ��2>@�����H�?             "@        I       J                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        N       O                 �n6@���Q��?	             $@        ������������������������       �                     @        P       U                     �?�q�q�?             @        Q       R                    �?�q�q�?             @        ������������������������       �                     �?        S       T                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        W       X                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        [       �                    �?��*���?E           �@       \       �                    �?Ȩ��?�            �x@        ]       x                 Ь*'@@�҇��?9            �W@        ^       u                    �?�\��N��?             C@       _       t                   �J@     ��?             @@       `       q                  �m#@X�Cc�?             <@       a       d                   �3@�\��N��?             3@        b       c                 P��@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        e       f                   �6@���Q��?             .@        ������������������������       �                     @        g       l                 P�@�eP*L��?             &@        h       k                   �9@      �?             @       i       j                    8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        m       n                 ��� @����X�?             @        ������������������������       �                     @        o       p                 `��!@      �?             @        ������������������������       �                      @        ������������������������       �                      @        r       s                 pF%@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        v       w                 P�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        y       �                    �?4և����?!             L@       z       �                     @$�q-�?             J@       {       �                   �*@��<D�m�?            �H@        |       }                 `f�)@"pc�
�?             &@        ������������������������       �                     �?        ~                          �B@z�G�z�?             $@       ������������������������       �                     @        �       �                    D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 `fF:@P�Lt�<�?             C@        �       �                     �?�}�+r��?
             3@        ������������������������       �                     @        �       �                    �?��S�ۿ?             .@        ������������������������       �                     @        �       �                   @B@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     3@        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �9@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     �?��$8�'�?�            �r@        �       �                   �<@p�ݯ��?$            �L@        �       �                 `f&F@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �>@�\�u��?             �I@        �       �                 ��$:@      �?             8@        ������������������������       �                     @        �       �                   @>@p�ݯ��?             3@       �       �                 03k:@��S���?	             .@        ������������������������       �                     @        �       �                   @=@�q�q�?             (@       �       �                 `f�;@�q�q�?             "@       �       �                   �K@և���X�?             @       �       �                 X��B@���Q��?             @        ������������������������       �                     �?        �       �                    H@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���R@PN��T'�?             ;@       ������������������������       �                     6@        �       �                  �6f@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �?�@��sK�z�?�            �n@        �       �                 P�N@@uvI��?>            �X@       ������������������������       �        $            �M@        �       �                 �Yu@ ���J��?            �C@        �       �                    �?      �?             @       �       �                    :@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �A@        �       �                 ��i @����?]            �b@        �       �                    �?r�q��?             H@       �       �                 @3�@"pc�
�?             F@        �       �                    �?z�G�z�?             $@       �       �                   �A@�����H�?             "@       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     �?        �       �                   �3@@�0�!��?             A@        �       �                   �2@�q�q�?             "@       �       �                    1@z�G�z�?             @       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     9@        ������������������������       �                     @        �       �                    �?P���Q�?@             Y@       �       �                   �@@(�s���?0             U@       �       �                     @0�)AU��?!            �L@        ������������������������       �                     7@        �       �                 @�!@г�wY;�?             A@        �       �                    8@�8��8��?             (@       ������������������������       �                     "@        �       �                   �=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        �       �                     @PN��T'�?             ;@       �       �                    F@8�Z$���?             :@        �       �                   @D@������?             .@       �       �                   �'@"pc�
�?             &@        ������������������������       �                     �?        �       �                   �A@z�G�z�?             $@        ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     0@        �       �                    �?�O
��?M            @]@        �       �                    B@b�h�d.�?            �A@       �       �                    �?(;L]n�?             >@       ������������������������       �        
             4@        �       �                 039@ףp=
�?             $@       �       �                 `f7@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @�=���D�?9            �T@        �       �                    @ҳ�wY;�?             1@       �       �                    �?ףp=
�?             $@       ������������������������       �                     @        �       �                 �(\�?�q�q�?             @        ������������������������       �                     �?        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @����X�?             @       �       �                 ���A@r�q��?             @        �       �                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �                       ���R@؇>���?,            @P@       �                           @�k�'7��?&            �L@        �                          �?�eP*L��?	             &@       �                         �L@���Q��?             $@       �                            �?      �?              @        ������������������������       �                      @                                 �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?                                 �?���}<S�?             G@                                @\-��p�?             =@             	                03c"@��s����?             5@        ������������������������       �                      @        
                      �|Y>@�KM�]�?             3@       ������������������������       �                     *@                                  @�q�q�?             @        ������������������������       �                     �?                                 @z�G�z�?             @        ������������������������       �                     @                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     1@                                 M@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub��������������"`c�?ȃ޺?9�?m����g�?&���0�?�=�����?��=���?��Moz��?Y�B��?      �?        ��.���?t�E]t�?              �?=��<���?�a�a�?              �?ffffff�?�������?      �?        �������?UUUUUU�?      �?              �?      �?�m۶m��?�$I�$I�?              �?�9�s��?�c�1��?]t�E]�?F]t�E�?�������?�������?      �?                      �?      �?        �������?�������?      �?      �?              �?      �?              �?        �&!����?�l�:��?�����?�ȍ�ȍ�?'�l��&�?6�d�M6�?Cy�5��?^Cy�5�?;�;��?;�;��?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?S�n0�?�Y7�"��?�4M�4M�?Y�eY�e�?ZLg1���?Lg1��t�?ڨ�l�w�?L� &W�?333333�?333333�?      �?      �?      �?        �������?�������?      �?      �?              �?      �?              �?              �?        h/�����?/�����?{�G�z�?
ףp=
�?      �?        �������?�������?              �?wwwwww�?�?      �?      �?              �?      �?        ]t�E�?F]t�E�?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?      �?                      �?�������?333333�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        UUUUUU�?�������?              �?      �?              �?        ����?�+�+�+�?w#-"�t�?�����?}g���Q�?!&W�+�?�5��P�?y�5���?      �?      �?�m۶m��?%I�$I��?�5��P�?y�5���?      �?      �?              �?      �?        �������?333333�?              �?t�E]t�?]t�E�?      �?      �?      �?      �?              �?      �?                      �?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?        �q�q�?�q�q�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        �m۶m۶?I�$I�$�?;�;��?�؉�؉�?և���X�?��S�r
�?F]t�E�?/�袋.�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?(�����?���k(�?(�����?�5��P�?              �?�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?DP/��M�?�}�>*��?^Cy�5�?Cy�5��?UUUUUU�?�������?              �?      �?        �������?�?      �?      �?      �?        Cy�5��?^Cy�5�?�������?�?              �?�������?�������?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?�������?333333�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?              �?&���^B�?h/�����?      �?        �������?�������?              �?      �?        .����-�?#6�a#�?�Cc}h��?9/���?      �?        ��-��-�?�A�A�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        S�n0�?�g�`�|�?�������?UUUUUU�?/�袋.�?F]t�E�?�������?�������?�q�q�?�q�q�?      �?              �?      �?              �?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?      �?      �?              �?        ffffff�?�������?�a�a�?��y��y�?��Gp�?p�}��?      �?        �?�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        &���^B�?h/�����?;�;��?;�;��?wwwwww�?�?/�袋.�?F]t�E�?      �?        �������?�������?�m۶m��?�$I�$I�?      �?              �?      �?      �?              �?              �?        �
��
��?���?_�_��?;��:���?�?�������?              �?�������?�������?      �?      �?              �?      �?                      �?      �?        w%jW�v�?�+Q��?�������?�������?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�m۶m��?�$I�$I�?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�����? �����?-����b�?Lg1��t�?]t�E�?t�E]t�?�������?333333�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ӛ���7�?d!Y�B�?a����?�{a���?z��y���?�a�a�?              �?�k(���?(�����?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?              �?      �?              �?              �?              �?      �?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJpVhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       d                    �?�C�"���?�           8�@                                   �?�F.< �?�            �p@                                    @��y� �?5            @W@        ������������������������       �                     G@                                   �?t/*�?            �G@                                   @������?             .@        ������������������������       �                     @                                   �?���Q��?             $@        	       
                 03�-@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                �|Y3@      �?             @        ������������������������       �                      @                                P�h2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                �|�9@      �?             @@        ������������������������       �                     $@                                   �?"pc�
�?             6@                                  �?������?
             .@                               ���@8�Z$���?	             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     @               U                    @�����?j            `e@                                   @NU��b��?Z            �a@        ������������������������       �        	             0@               $                 `f�$@@�j���?Q            @_@                                  �3@���|���?             6@        ������������������������       �                     @                #                  sW@@�0�!��?             1@        !       "                   �@@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        %       J                    �?�v�G���?D            �Y@       &       =                   �E@ףp=
�?5             T@       '       <                   �?@����?*            @P@       (       1                     @��-�=��?            �C@       )       *                     �?�g�y��?             ?@        ������������������������       �                     (@        +       0                    �?�}�+r��?
             3@       ,       -                    �?$�q-�?             *@       ������������������������       �                     @        .       /                   �7@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        2       3                    �?      �?              @        ������������������������       �                      @        4       ;                 `fV6@      �?             @       5       :                    �?���Q��?             @       6       9                 ��1@      �?             @       7       8                 �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        >       ?                   @F@������?             .@        ������������������������       �                      @        @       I                    �?8�Z$���?
             *@       A       B                    G@r�q��?	             (@        ������������������������       �                     @        C       H                     @�<ݚ�?             "@       D       G                   �*@      �?              @        E       F                   �J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        K       L                    ,@�û��|�?             7@        ������������������������       �                     @        M       N                     @�z�G��?             4@       ������������������������       �                     (@        O       P                 @34@      �?              @        ������������������������       �                     �?        Q       R                    @؇���X�?             @       ������������������������       �                     @        S       T                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        V       c                    @�������?             >@       W       `                 �|�:@�X����?             6@       X       Y                      @��
ц��?	             *@        ������������������������       �                      @        Z       [                   -@���|���?             &@        ������������������������       �                     @        \       ]                    �?      �?              @        ������������������������       �                      @        ^       _                 ��T?@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        a       b                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        e       �                    �?��H�&p�?           �{@        f       �                 ��<J@.�	F�9�?3            @T@       g       p                     @PN��T'�?$             K@        h       o                     �?�C��2(�?             6@       i       n                  Y>@r�q��?	             (@        j       k                 ���<@      �?             @        ������������������������       �                     �?        l       m                 X��E@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        q       �                 03�-@     ��?             @@       r       w                   �5@؇���X�?             <@        s       t                    �?�q�q�?             @        ������������������������       �                     �?        u       v                    -@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        x       �                    �?HP�s��?             9@       y       �                 �|�=@�C��2(�?             6@       z                          @@�r����?
             .@       {       |                 ���@�8��8��?             (@        ������������������������       �                     @        }       ~                 �|=@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        �       �                 ��� @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�q�q�?             ;@       �       �                  �}S@      �?             0@        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        ������������������������       �                     @        �       �                   �H@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�C��2(�?             &@       ������������������������       �                     @        �       �                 �\@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    #@r�q��?�            �v@        �       �                 @3�4@��}*_��?             ;@        ������������������������       �                     $@        �       �                    �?j���� �?
             1@        ������������������������       �                     �?        �       �                    @     ��?	             0@        ������������������������       �                     @        ������������������������       �                     "@        �       �                     �?�����?�            0u@        �       �                    �?�q�q�?$            �O@       �       �                    �?��Q��?!             N@       �       �                 �|�<@�q�q�?             H@        �       �                 `f�D@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @E@���?            �D@        ������������������������       �                     0@        �       �                    @@���Q��?             9@       �       �                    L@�\��N��?
             3@       �       �                   `G@      �?             (@        �       �                   �F@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    R@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                  x#J@�q�q�?             (@        ������������������������       �                     @        �       �                   �B@X�<ݚ�?             "@       �       �                    <@�q�q�?             @        ������������������������       �                     �?        �       �                    >@z�G�z�?             @        ������������������������       �                     @        �       �                 `f�K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�8��8��?�            @q@       �       �                 �?�@�W�l~�?�             l@        �       �                    �?�nkK�?>             W@        �       �                 ��(@�KM�]�?             3@       �       �                 ���@      �?             0@        ������������������������       �                      @        �       �                 �|Y=@؇���X�?	             ,@        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     @        �       �                 ���@��pBI�?2            @R@        �       �                 ���@��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        �       �                    ?@ _�@�Y�?(             M@       ������������������������       �        !            �G@        �       �                   @@@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?؇���X�?V            �`@        ������������������������       �                      @        �       �                     @�������?U            ``@        �       �                   �*@�L���?            �B@       �       �                    5@ףp=
�?             >@        �       �                    &@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|Y=@�>����?             ;@        ������������������������       �                     (@        �       �                 `f�)@�r����?             .@        ������������������������       �                     @        �       �                 �|�=@"pc�
�?             &@        ������������������������       �                     �?        �       �                   �C@ףp=
�?             $@        ������������������������       �                     @        �       �                    G@؇���X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �;@t/*�?8            �W@        �       �                    9@��X��?             <@       �       �                 0S5 @�q�q�?             8@        �       �                   �3@�eP*L��?             &@        �       �                   �2@����X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �        
             *@        ������������������������       �                     @        �       �                   �>@��IF�E�?$            �P@        �       �                 `��!@������?             B@       �       �                 �|Y=@      �?
             0@        ������������������������       �                     @        �       �                 �|�=@$�q-�?	             *@       �       �                 ��) @�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        �       �                 @3�@z�G�z�?             >@        �       �                   �A@���Q��?             $@       �       �                   �?@�q�q�?             "@        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �        #            �I@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������[�e�?���I54�?>����?|��|�?X`��??���O?�?              �?W�+���?�;����?�?wwwwww�?              �?�������?333333�?      �?      �?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?      �?      �?              �?F]t�E�?/�袋.�?�?wwwwww�?;�;��?;�;��?      �?                      �?      �?                      �?^Cy�5�?Q^Cy��?qJ��O$�?d-C���?              �?X9��v��?���Mb�?]t�E]�?F]t�E�?              �?ZZZZZZ�?�������?      �?      �?              �?      �?              �?        ��O �?C���?�������?�������? �����?~�~��?�A�A�?}˷|˷�?�B!��?��{���?              �?(�����?�5��P�?;�;��?�؉�؉�?              �?UUUUUU�?�������?      �?                      �?              �?      �?      �?              �?      �?      �?�������?333333�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?                      �?�?wwwwww�?      �?        ;�;��?;�;��?UUUUUU�?�������?              �?�q�q�?9��8���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?��,d!�?8��Moz�?      �?        333333�?ffffff�?              �?      �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        �������?�������?�E]t��?]t�E]�?�;�;�?�؉�؉�?              �?]t�E]�?F]t�E�?              �?      �?      �?      �?        �������?UUUUUU�?      �?                      �?�q�q�?�q�q�?              �?      �?              �?        ��o�j�?�IA��U�?�����H�?~X�<��?&���^B�?h/�����?]t�E�?F]t�E�?�������?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        q=
ףp�?{�G�z�?]t�E�?F]t�E�?�������?�?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?�������?�������?      �?              �?      �?              �?      �?        ]t�E�?F]t�E�?      �?        �������?�������?              �?      �?        �������?UUUUUU�?B{	�%��?_B{	�%�?              �?�������?ZZZZZZ�?      �?              �?      �?              �?      �?        ���G���?.�	���?UUUUUU�?UUUUUU�?�������?ffffff�?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?      �?        28��1�?8��18�?      �?        333333�?�������?�5��P�?y�5���?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?      �?        �������?�������?      �?        �q�q�?r�q��?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?2Tv���?�o^M<+�?�Mozӛ�?d!Y�B�?�k(���?(�����?      �?      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?        ���Ǐ�?����?�������?�?      �?                      �?#,�4�r�?�{a���?      �?        ]t�E�?F]t�E�?              �?      �?        ۶m۶m�?�$I�$I�?      �?        #����[�?s�U���?}���g�?L�Ϻ��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?        �Kh/��?h/�����?      �?        �������?�?      �?        /�袋.�?F]t�E�?              �?�������?�������?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?        �;����?W�+���?n۶m۶�?%I�$I��?UUUUUU�?�������?t�E]t�?]t�E�?�$I�$I�?�m۶m��?              �?      �?      �?      �?              �?                      �?�l��&��?'�l��&�?�q�q�?�q�q�?      �?      �?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM+hjh))��}�(h,h/h0M+��h2h3h4hph<�h=Kub������       n                 ���$@���$ӡ�?�           8�@                                  �0@���ۜ1�?�            �p@                                   �?      �?              @       ������������������������       �                     @                                pf�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                �ٝ@f?�ϼ��?�            `p@        	       
                 ���@����Q8�?)            �Q@        ������������������������       �                    �@@                                   7@�KM�]�?             C@        ������������������������       �                     @                                   �?      �?             @@                               ���@@�0�!��?             1@                               X��B@z�G�z�?             $@                               �|Y;@      �?              @        ������������������������       �                     �?                                   �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                �|�=@؇���X�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                      @                                ���@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@               #                    �?P/�DGT�?t            �g@                                �|Y=@<=�,S��?            �A@        ������������������������       �                     @               "                    �?     ��?             @@                !                    �?�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     5@        $       1                   �2@���B���?_            �c@        %       &                   �1@�n_Y�K�?             *@        ������������������������       �                     �?        '       .                    �?�q�q�?             (@       (       -                    �?և���X�?             @       )       *                 P��@�q�q�?             @        ������������������������       �                     @        +       ,                 ��!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        /       0                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        2       ]                 �|�=@$���'w�?X            �a@       3       D                    �?t�6Z���?B            �[@        4       A                    �?և���X�?
             ,@       5       @                    ;@�q�q�?             (@       6       7                   �4@�z�G��?             $@        ������������������������       �                     �?        8       ?                 03�!@�<ݚ�?             "@       9       :                 ���@      �?              @        ������������������������       �                     @        ;       >                   �9@      �?             @       <       =                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        B       C                 �!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        E       F                 �?�@�8��8��?8             X@        ������������������������       �                     H@        G       \                 �|Y=@r�q��?             H@       H       S                   �:@�<ݚ�?             B@       I       R                   �4@8�Z$���?             :@       J       Q                    �?      �?	             0@       K       P                 0S5 @z�G�z�?             .@        L       M                 @3�@�q�q�?             "@        ������������������������       �                      @        N       O                   �3@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        T       [                    �?���Q��?             $@       U       V                 0S%"@և���X�?             @        ������������������������       �                     @        W       X                   �<@      �?             @        ������������������������       �                      @        Y       Z                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ^       g                   @@@���!pc�?            �@@        _       b                   �>@��
ц��?	             *@        `       a                 �̌!@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        c       d                 P�@�q�q�?             "@        ������������������������       �                      @        e       f                   �?@և���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        h       i                   �B@ףp=
�?             4@       ������������������������       �                     "@        j       k                    �?"pc�
�?             &@        ������������������������       �                     �?        l       m                   �C@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        o       �                  x#J@�k����?           �{@       p       y                    @� ���?�            Pt@        q       r                    @���j��?             G@       ������������������������       �                     @@        s       t                 ��T?@@4և���?	             ,@       ������������������������       �                     "@        u       x                    @z�G�z�?             @       v       w                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        z       �                   �K@pY���?�            pq@       {       �                    �?�K)��;�?�            �p@        |       }                   �-@��U/��?L            �\@        ������������������������       �                     @        ~       �                     @ҷ{�&�?G            �Z@              �                 `f�)@����?*            @P@        ������������������������       �                     (@        �       �                    �?�NW���?"            �J@       �       �                   �B@$�q-�?!             J@       �       �                    �?г�wY;�?             A@       �       �                    �?P���Q�?             4@        ������������������������       �                     @        �       �                   �7@��S�ۿ?
             .@        �       �                    ?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �        	             ,@        �       �                    �?r�q��?
             2@        �       �                    �?�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @F@�����H�?             "@        �       �                   �E@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��p@@��6���?             E@       �       �                 ��T?@�ʻ����?             A@       �       �                    �?     ��?             @@       �       �                    �?�g�y��?             ?@        �       �                    �?�q�q�?
             .@        �       �                 ���,@      �?              @        ������������������������       �                     @        �       �                  S�-@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03�-@և���X�?             @        ������������������������       �                     @        �       �                 `�@1@      �?             @       �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �B@      �?             0@       �       �                    �?��
ц��?             *@       �       �                 `fV6@�q�q�?
             (@       �       �                    �?      �?	             $@       �       �                 �|�;@      �?              @        ������������������������       �                     @        �       �                   �>@z�G�z�?             @        ������������������������       �                      @        �       �                 03�1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 `fv1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?B�`�?^            �b@       �       �                 ��$:@Ȩ�I��??            �Z@       �       �                     @ 	��p�?$             M@       �       �                    �?`'�J�?            �I@        ������������������������       �                     @        �       �                    5@`�q�0ܴ?            �G@        �       �                   �'@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �C@ qP��B�?            �E@       ������������������������       �                     :@        �       �                    ,@�IєX�?
             1@       �       �                   �F@      �?              @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     "@        �       �                 ��q1@����X�?             @       ������������������������       �                     @        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             H@        �       �                 `f�A@���Q��?             $@       �       �                  �>@և���X�?             @       �       �                  Y>@���Q��?             @       �       �                 �|�=@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �G@�\��N��?             C@       �       �                    G@�f7�z�?             =@       �       �                 ��yC@��
ц��?             :@       �       �                    D@z�G�z�?	             .@       �       �                 �|�<@�8��8��?             (@        ������������������������       �                     @        �       �                   `@@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     &@        ������������������������       �                     @        �       �                   �J@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                    $@�:�^���?            �F@        �       �                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �5@������?            �D@        �       �                    �?r�q��?             @       �       �                    2@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @��?^�k�?            �A@        ������������������������       �                     *@        �       �                 ��.@���7�?             6@        �       �                    �?      �?             @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             2@        ������������������������       �                     ,@        �       *                  �O@�c�Α�?I             ]@              %                `fmj@x��}�?F            �[@             "                   F@��!���?<            @W@                                 �?�ӖF2��?-            �Q@                                �?�����H�?'            �O@                                �?�(\����?             D@       ������������������������       �                     C@                                �0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        	                         �?��+7��?             7@       
                        �8@���|���?             &@                             ���Q@�q�q�?             @        ������������������������       �                     �?                                 �?z�G�z�?             @                               �4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 �?r�q��?             (@                               �B@      �?              @                             ���M@�q�q�?             @                                @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 ;@      �?              @                                 �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?               !                �|�>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        #      $                   �?���|���?             6@       ������������������������       �        	             ,@        ������������������������       �                      @        &      )                X�,@@j���� �?
             1@       '      (                `f�n@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M+KK��h2h3h4hVh<�h=Kub������������H�1�N�?oݟ�Kb�?�b���?�u�< �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�]�WqB�?ˈ>�:��?O�o�z2�?��Vج?      �?        �k(���?(�����?      �?              �?      �?ZZZZZZ�?�������?�������?�������?      �?      �?      �?        �m۶m��?�$I�$I�?              �?      �?              �?        ۶m۶m�?�$I�$I�?�������?�������?      �?        �������?�?              �?      �?        ���M���?���?�A�A�?X|�W|��?              �?      �?      �?F]t�E�?]t�E�?              �?      �?              �?        ��؉���?ى�؉��?;�;��?ى�؉��?      �?        �������?�������?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?              �?      �?        �w��g�?9 2ܫ`�?X���oX�?��)A��?۶m۶m�?�$I�$I�?�������?�������?333333�?ffffff�?      �?        �q�q�?9��8���?      �?      �?              �?      �?      �?      �?      �?              �?      �?                      �?      �?              �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?9��8���?�q�q�?;�;��?;�;��?      �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?              �?                      �?      �?        333333�?�������?۶m۶m�?�$I�$I�?              �?      �?      �?      �?              �?      �?      �?                      �?      �?              �?        F]t�E�?t�E]t�?�؉�؉�?�;�;�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?              �?      �?      �?�������?�������?      �?        /�袋.�?F]t�E�?      �?        �������?�������?              �?      �?        ���g5��?'�L��?�����?�ȍ�ȍ�?!Y�B�?ozӛ���?              �?n۶m۶�?�$I�$I�?      �?        �������?�������?      �?      �?      �?                      �?      �?        ҝ̇t'�?\�f���?ߑa��y�?B�<���?g1��t�?Lg1��t�?      �?        !V��G&�?�Ե���? �����?~�~��?              �?�x+�R�?萚`���?;�;��?�؉�؉�?�?�?�������?ffffff�?              �?�?�������?      �?      �?      �?                      �?              �?              �?UUUUUU�?�������?�q�q�?9��8���?      �?              �?      �?      �?                      �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?              �?b�a��?=��<���?<<<<<<�?�������?      �?      �?��{���?�B!��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?�;�;�?�؉�؉�?�������?�������?      �?      �?      �?      �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?      �?                      �?      �?                      �?              �?      �?        ���o�7�?ـl@6 �?+�R��?�	�[���?������?�{a���?�������?�?      �?        ��F}g��?W�+�ɥ?      �?      �?              �?      �?        ��}A�?�}A_З?      �?        �?�?      �?      �?      �?      �?      �?              �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?333333�?�������?۶m۶m�?�$I�$I�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �5��P�?y�5���?O#,�4��?a���{�?�;�;�?�؉�؉�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?        �q�q�?�q�q�?              �?      �?        }�'}�'�?l�l��?      �?      �?              �?      �?        p>�cp�?������?�������?UUUUUU�?�������?�������?      �?                      �?      �?        _�_��?�A�A�?      �?        �.�袋�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        �{a���?5�rO#,�?A��)A�?pX���o�?'�h��&�?v�e�]v�?�z2~���?Zas �
�?�q�q�?�q�q�?�������?333333�?              �?      �?      �?      �?                      �?Y�B��?zӛ����?F]t�E�?]t�E]�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?              �?      �?              �?                      �?UUUUUU�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?              �?      �?      �?      �?      �?              �?      �?              �?      �?      �?                      �?F]t�E�?]t�E]�?              �?      �?        ZZZZZZ�?�������?ffffff�?333333�?      �?                      �?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��nhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������                           @�,�٧��?�           8�@               	                    �?�'�`d�?            �@@                                 �C@�J�4�?             9@                                  �?���}<S�?             7@       ������������������������       �                     *@                                   @z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        
                           @      �?              @                                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                  @:HJ���?�           0�@              �                    �?��œ�L�?�           x�@              6                    �?����?S           ��@               !                    �?\X��t�?V            @a@                                  �-@p��%���?'            @Q@                                   �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                                ���@      �?%             P@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �E@0�z��?�?#             O@       ������������������������       �                     L@                                    �?r�q��?             @                                ,w�U@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        "       )                 �|Y<@��X���?/            @Q@        #       $                    3@����X�?	             ,@        ������������������������       �                     �?        %       (                 ���0@�θ�?             *@       &       '                   �6@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        *       5                 p�w@�1�`jg�?&            �K@       +       4                    �?�O4R���?%            �J@       ,       3                     �?h�����?             <@        -       2                 �|�=@ףp=
�?	             $@        .       1                 ��2>@      �?             @        /       0                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     9@        ������������������������       �                      @        7       �                    �?�X�~�?�            �x@       8       O                    �?fv�S��?�            �t@        9       :                   �5@X�;�^o�?#            �K@        ������������������������       �                     $@        ;       @                   �9@���V��?            �F@        <       ?                 pff@���|���?             &@        =       >                    8@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        A       B                 �Y5@l��\��?             A@        ������������������������       �                     �?        C       F                 ��� @�FVQ&�?            �@@        D       E                 �|�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        G       H                     �?(;L]n�?             >@        ������������������������       �                     &@        I       N                     @�}�+r��?             3@       J       M                   �*@�X�<ݺ?             2@       K       L                   �B@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        P       �                   @S@��-�=��?�            q@       Q       v                 �|�=@|0M�Y4�?�            �p@       R       Y                     �? eD5�Ҽ?k            �d@        S       T                 �|Y=@R���Q�?             4@        ������������������������       �                      @        U       V                 `fF<@r�q��?
             2@        ������������������������       �                     "@        W       X                   �>@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        Z       _                     @���N8�?`            `b@        [       ^                    4@      �?             @@        \       ]                    &@�8��8��?             (@        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                     4@        `       u                 �|Y=@P���Q�?N            �\@       a       l                 ���"@p��@���?:            @U@       b       e                 ���@��?^�k�?1            �Q@        c       d                 ���@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        f       g                 @3�@0�z��?�?+             O@       ������������������������       �                    �E@        h       k                   �2@�}�+r��?             3@        i       j                 ��Y @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             ,@        m       p                 `�X#@������?	             .@        n       o                   �8@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        q       r                 �!&B@�C��2(�?             &@       ������������������������       �                      @        s       t                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     >@        w       �                     �?8�Z$���?A             Z@        x       �                   �J@`�Q��?             9@       y       �                   �G@D�n�3�?             3@       z       {                 ��:@     ��?	             0@        ������������������������       �                     @        |                          �F@      �?             $@       }       ~                   @@@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                     @$��$�L�?0            �S@        �       �                   �*@�����H�?             ;@       �       �                   �C@@�0�!��?             1@        ������������������������       �                     @        �       �                   �F@�z�G��?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     $@        �       �                   @@@4��?�?              J@        �       �                 �̌!@�z�G��?             $@       �       �                    ?@      �?              @        ������������������������       �                     @        �       �                   �@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@���N8�?             E@       ������������������������       �                     4@        �       �                 @3�@�C��2(�?             6@        ������������������������       ��q�q�?             @        ������������������������       �        
             3@        ������������������������       �                      @        �       �                 039@
;&����?-            @Q@        �       �                    �?������?             ;@       �       �                     @��
ц��?	             *@        ������������������������       �                     �?        �       �                 �|�;@      �?             (@        �       �                    6@r�q��?             @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���.@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    6@@4և���?             ,@        �       �                    3@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     �?�ՙ/�?             E@       �       �                   �I@J�8���?             =@       �       �                    �?���Q��?             9@       �       �                    �?�q�q�?             8@        ������������������������       �                      @        �       �                  x#J@      �?
             0@        ������������������������       �                     @        �       �                   @K@      �?             (@        ������������������������       �                     @        �       �                   �D@      �?              @        �       �                 `f�N@�q�q�?             @        ������������������������       �                     �?        �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �:@��
ц��?
             *@        ������������������������       �                      @        �       �                    �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                    D@r�q��?P             ^@       �       �                    @@��Pl3�?C            @X@       �       �                     @\Ќ=��??            �V@       �       �                   �(@���c�H�?$            �H@        ������������������������       �                      @        �       �                    �?��k=.��?#            �G@        �       �                    �?և���X�?             ,@        ������������������������       �                     @        �       �                    �?      �?              @       �       �                    �?z�G�z�?             @       �       �                    >@      �?             @        ������������������������       �                      @        �       �                 �;�p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                  "&d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�C��2(�?            �@@       ������������������������       �                     >@        ������������������������       �                     @        �       �                    3@�D����?             E@        �       �                 ���4@      �?             4@       �       �                  S%/@�n_Y�K�?             *@       �       �                    �?      �?              @       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    +@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `v�6@�eP*L��?             6@       �       �                 �=/@�q�q�?             2@       �       �                 �|�?@�eP*L��?             &@       �       �                    �?      �?              @       �       �                 �|�<@      �?             @        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                     @r�q��?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                 ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �                           @��<b���?             7@       �                          @I@�t����?
             1@        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                  �?r�q��?             (@                               �K@�C��2(�?             &@        ������������������������       �                     @                                 �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        	                         @�nkK�?             7@       
                      hf�2@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     (@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������&��jq�?:�g *�?'�l��&�?6�d�M6�?{�G�z�?�z�G��?d!Y�B�?ӛ���7�?              �?�������?�������?              �?      �?              �?              �?      �?333333�?�������?              �?      �?                      �?��@n�?�~#���?=\��D��?�G�lv��?j�Ǡ��?-U�q�^�?��Moz��?!Y�B�?ہ�v`��?�g��%�?�������?333333�?              �?      �?              �?      �?      �?      �?              �?      �?        �B!��?|���{�?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?�Q�g���?��v`��?�$I�$I�?�m۶m��?      �?        �؉�؉�?ى�؉��?۶m۶m�?�$I�$I�?              �?      �?                      �?A��)A�?�־a�?:�&oe�?�x+�R�?�m۶m��?�$I�$I�?�������?�������?      �?      �?      �?      �?      �?                      �?      �?              �?              �?              �?                      �?s�$��6�?}��`��?��]�ڕ�?�]�ڕ��?J��yJ�?�־a��?              �?�>�>��?[�[��?F]t�E�?]t�E]�?      �?      �?              �?      �?              �?        �������?------�?      �?        |���?>����?UUUUUU�?UUUUUU�?              �?      �?        �?�������?              �?(�����?�5��P�?�q�q�?��8��8�?�������?�������?              �?      �?                      �?              �?}˷|˷�?�A�A�?P��9��?~�3���?:�2	v�?\��l���?333333�?333333�?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��y��y�?�a�a�?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        �ø_�T�?��s���?�������?�?_�_��?�A�A�?      �?      �?      �?                      �?|���{�?�B!��?      �?        �5��P�?(�����?�������?�������?              �?      �?              �?        wwwwww�?�?      �?      �?      �?                      �?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ;�;��?;�;��?��(\���?{�G�z�?l(�����?(������?      �?      �?      �?              �?      �?�$I�$I�?�m۶m��?      �?                      �?      �?                      �?      �?        ��]-n��?�3���?�q�q�?�q�q�?ZZZZZZ�?�������?      �?        ffffff�?333333�?      �?      �?      �?              �?        �N��N��?ى�؉��?ffffff�?333333�?      �?      �?      �?        �������?�������?              �?      �?                      �?��y��y�?�a�a�?      �?        ]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?Y�B��?�Mozӛ�?B{	�%��?{	�%���?�;�;�?�؉�؉�?      �?              �?      �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        UUUUUU�?�������?      �?                      �?n۶m۶�?�$I�$I�?�������?UUUUUU�?      �?                      �?      �?        �a�a�?�<��<��?|a���?�rO#,��?�������?333333�?�������?�������?              �?      �?      �?      �?              �?      �?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?              �?�؉�؉�?�;�;�?      �?        F]t�E�?]t�E]�?              �?      �?        UUUUUU�?UUUUUU�?�n�'�i�?��4l7��?�Q�Q�?s5Ws5W�?/�����?4և����?      �?        br1���?g���Q��?۶m۶m�?�$I�$I�?              �?      �?      �?�������?�������?      �?      �?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        F]t�E�?]t�E�?              �?      �?        �0�0�?z��y���?      �?      �?;�;��?ى�؉��?      �?      �?      �?              �?      �?              �?      �?        �������?�������?              �?      �?              �?        ]t�E�?t�E]t�?UUUUUU�?UUUUUU�?t�E]t�?]t�E�?      �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?              �?      �?              �?                      �?      �?        UUUUUU�?�������?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?��,d!�?��Moz��?�������?�������?�������?333333�?              �?      �?        �������?UUUUUU�?]t�E�?F]t�E�?      �?        �������?�������?              �?      �?                      �?      �?        �Mozӛ�?d!Y�B�?]t�E�?F]t�E�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJXk�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM'hjh))��}�(h,h/h0M'��h2h3h4hph<�h=Kub������       x                     @�,�٧��?�           8�@                                  �2@F���V�?�            �t@        ������������������������       �                    �@@               K                     �?�����?�            �r@              @                    �?J�8���?c            �e@                                  �?�9!���?Q            �a@               
                 03�=@@3����?             K@               	                   �H@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �I@               ;                   �H@ƈ�VM�?2            @V@                                  �?�;�vv��?'            @R@                                X�,@@�	j*D�?
             :@                               0��G@�q�q�?             (@                                 Y>@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                �|Y;@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@                                ��I/@֭��F?�?            �G@        ������������������������       �                     @               *                   �>@�>$�*��?            �D@               )                   @>@p�ݯ��?             3@                               03k:@      �?	             ,@        ������������������������       �                     �?                                  �<@��
ц��?             *@        ������������������������       �                     �?                                 �|Y=@�q�q�?             (@        ������������������������       �                      @        !       (                   @=@      �?             $@       "       #                 �|�?@      �?              @        ������������������������       �                      @        $       %                   �C@      �?             @        ������������������������       �                      @        &       '                 `f�;@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        +       0                    �?���!pc�?             6@        ,       -                   �A@�����H�?             "@        ������������������������       �                     @        .       /                 ��yC@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        1       :                    �?�n_Y�K�?             *@       2       9                 03�U@�q�q�?             (@       3       8                 ���L@�<ݚ�?             "@        4       5                    7@      �?             @        ������������������������       �                     �?        6       7                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        <       ?                    �?      �?             0@       =       >                   �R@$�q-�?
             *@       ������������������������       �        	             (@        ������������������������       �                     �?        ������������������������       �                     @        A       J                   �L@��a�n`�?             ?@       B       I                    �?؇���X�?             <@        C       D                 03/O@�q�q�?             (@        ������������������������       �                     @        E       F                    �?�����H�?             "@       ������������������������       �                     @        G       H                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     @        L       q                    �?b �y��?P            �_@       M       X                   �(@">�֕�?@            @Z@        N       Q                   �@@�J�4�?             9@       O       P                    5@P���Q�?             4@        ������������������������       ��q�q�?             @        ������������������������       �        
             1@        R       S                   @A@���Q��?             @        ������������������������       �                      @        T       U                   @E@�q�q�?             @        ������������������������       �                     �?        V       W                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Y       d                    �?�G�z��?0             T@        Z       a                   �B@r�q��?             >@       [       `                   �7@ȵHPS!�?             :@       \       ]                    �?@�0�!��?             1@        ������������������������       �                     @        ^       _                   �;@d}h���?
             ,@        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     "@        b       c                   �C@      �?             @        ������������������������       �                      @        ������������������������       �                      @        e       f                    �?HP�s��?             I@        ������������������������       �                     @        g       p                   �*@�C��2(�?             F@        h       m                   �C@"pc�
�?             6@       i       j                 �|Y;@��S�ۿ?	             .@        ������������������������       �                     @        k       l                 �|�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        n       o                   �F@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     6@        r       w                 ��J@      �?             6@       s       v                    �?�G�z��?             4@       t       u                    �?D�n�3�?             3@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                      @        y       &                   @0tE`��?�            �w@       z       �                  �#@�_q��>�?�            w@       {       |                 ���@ �y63��?�            �n@        ������������������������       �                     9@        }       �                    �?���z��?�            �k@        ~       �                   �3@8�$�>�?            �E@               �                    1@$�q-�?             *@        ������������������������       �                      @        �       �                   �2@z�G�z�?             @        �       �                 P��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �4@��S���?             >@        ������������������������       �                     @        �       �                    �?�5��?             ;@       �       �                  S�"@�q�q�?             8@       �       �                 ���@8����?             7@        ������������������������       �                      @        �       �                    �?�q�q�?             5@        �       �                 ���@z�G�z�?             $@        ������������������������       �                     �?        �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �6@�eP*L��?             &@        ������������������������       �                     @        �       �                 ��� @����X�?             @       �       �                    8@r�q��?             @        �       �                 @3�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                ��k @N�hƇ�?u             f@        ������������������������       �                     �?        �       �                    �?h�V���?t             f@       �       �                    �?���W���?p            �e@        �       �                   �6@�:�]��?            �I@        ������������������������       �                      @        �       �                    �?@9G��?            �H@       �       �                 �|Y?@(;L]n�?             >@       �       �                 �|=@���N8�?             5@        ������������������������       �                     @        �       �                 ���@�IєX�?
             1@        ������������������������       �                     @        �       �                   @@�C��2(�?             &@       ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     "@        �       �                  ��@�}�+r��?             3@        ������������������������       �                     @        �       �                 ��(@$�q-�?             *@       �       �                 �|Y=@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        �       �                 ���@����W1�?T            @^@        ������������������������       �                      @        �       �                 �?�@�D�d@6�?S            �]@        �       �                 �?$@�O4R���?'            �J@        �       �                 �|Y>@ �q�q�?             8@       �       �                 �|�;@�C��2(�?	             &@       ������������������������       �                      @        �       �                 ��,@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     =@        �       �                 �|�=@r�q��?,            �P@       �       �                   �3@�8��8��?              H@        �       �                 0S5 @�<ݚ�?             "@        �       �                   �1@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �:@�7��?            �C@        ������������������������       �                     1@        �       �                 ��) @�C��2(�?             6@       ������������������������       �                     *@        �       �                   �;@�<ݚ�?             "@        ������������������������       �                     �?        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �?@b�2�tk�?             2@        �       �                   �>@      �?             @       �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �F@����X�?	             ,@       �       �                 ��I @���|���?             &@       �       �                   �A@և���X�?             @       ������������������������       ��q�q�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?����-T�?M             _@        �       �                     @<=�,S��?            �A@       �       �                 X��B@����e��?            �@@       �       �                 03�7@f���M�?             ?@       �       �                    �?������?             ;@        �       �                 P��+@և���X�?             @        ������������������������       �                     @        �       �                 �0@      �?             @        ������������������������       �                      @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?z�G�z�?             4@       �       �                   �-@r�q��?             (@       �       �                    �?����X�?             @        �       �                   �,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?              @       �       �                 �|�4@r�q��?             @        ������������������������       �                      @        �       �                 ��.@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                               0S�*@���*~�?6            @V@                                �7@r�q��?             @       ������������������������       �                     @                                �=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 @4�{Y���?0            �T@              
                   �?���Q��?             $@              	                ��1<@      �?             @       ������������������������       �                      @        ������������������������       �                      @                                 @�q�q�?             @                                �?���Q��?             @        ������������������������       �                      @                              ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                 �?d1<+�C�?)            @R@                              pff0@�n_Y�K�?             *@        ������������������������       �                     @                              `fV6@r�q��?             @        ������������������������       �                     @                              �T)D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @              %                   �?�8��8��?!             N@                                 �?��hJ,�?             A@                              ��1@�	j*D�?             *@                              �|�;@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        !      $                   0@���N8�?             5@        "      #                  �/@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             0@        ������������������������       �                     :@        ������������������������       �                      @        �*       h�h))��}�(h,h/h0M'KK��h2h3h4hVh<�h=Kub�������������&��jq�?:�g *�?����f�?����L�?              �?�W���g�?3T1���?|a���?�rO#,��?̒r@d��?�����#�?h/�����?���Kh�?UUUUUU�?UUUUUU�?              �?      �?                      �?+Y�JV��?�MmjS��?�8�?����Ǐ�?;�;��?vb'vb'�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?        �������?333333�?              �?      �?                      �?�F}g���?br1���?      �?        �18���?�����?Cy�5��?^Cy�5�?      �?      �?              �?�;�;�?�؉�؉�?              �?�������?�������?      �?              �?      �?      �?      �?      �?              �?      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?        �������?�������?              �?      �?        ;�;��?ى�؉��?�������?�������?9��8���?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?              �?      �?�؉�؉�?;�;��?      �?                      �?      �?        �s�9��?�c�1��?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        :�N����?��b�X,�?_�_��?�A�A�?�z�G��?{�G�z�?ffffff�?�������?UUUUUU�?UUUUUU�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ffffff�?333333�?UUUUUU�?�������?�؉�؉�?��N��N�?�������?ZZZZZZ�?              �?۶m۶m�?I�$I�$�?      �?                      �?              �?      �?      �?      �?                      �?q=
ףp�?{�G�z�?      �?        ]t�E�?F]t�E�?/�袋.�?F]t�E�?�������?�?      �?              �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?              �?      �?�������?�������?l(�����?(������?              �?      �?                      �?              �?�A�χ�?�������?�M�0Z^�?1ɾ=���?0J5y��?�?�*��?      �?        *A��)�?X���oX�?�5eMYS�?6eMYS��?;�;��?�؉�؉�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�?      �?        /�����?h/�����?UUUUUU�?UUUUUU�?8��Moz�?d!Y�B�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?        �q�q�?�q�q�?              �?      �?        ]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?              �?        �z����?($�z�?              �?�袋.��?/�袋.�?*kʚ���?���)kʺ?}}}}}}�?�?              �?������?9/���?�������?�?��y��y�?�a�a�?      �?        �?�?      �?        ]t�E�?F]t�E�?�������?�������?      �?              �?        �5��P�?(�����?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?        ��eP*L�?���|���?              �?}��|���?���й?:�&oe�?�x+�R�?�������?UUUUUU�?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?9��8���?�q�q�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        ��[��[�?�A�A�?      �?        ]t�E�?F]t�E�?      �?        9��8���?�q�q�?              �?      �?      �?              �?      �?        �8��8��?9��8���?      �?      �?      �?      �?      �?                      �?              �?�m۶m��?�$I�$I�?]t�E]�?F]t�E�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?      �?              �?              �?        k���Zk�?)��RJ)�?X|�W|��?�A�A�?6�d�M6�?e�M6�d�?��Zk���?��RJ)��?{	�%���?B{	�%��?۶m۶m�?�$I�$I�?              �?      �?      �?      �?              �?      �?      �?                      �?�������?�������?UUUUUU�?�������?�$I�$I�?�m۶m��?      �?      �?              �?      �?        �������?�������?      �?                      �?              �?      �?      �?UUUUUU�?�������?              �?      �?      �?              �?      �?              �?      �?      �?                      �?      �?              �?                      �?���d%+�?��MmjS�?UUUUUU�?�������?              �?      �?      �?      �?                      �?�b��7��?4u~�!��?333333�?�������?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ݹs�Ν�?�1bĈ�?;�;��?ى�؉��?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?KKKKKK�?�������?vb'vb'�?;�;��?۶m۶m�?�$I�$I�?      �?                      �?      �?        ��y��y�?�a�a�?�������?�������?      �?                      �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ0��JhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       b                     @ʻ�J��?�           8�@                                  �1@���Ua��?�            t@        ������������������������       �                     :@                                   �?�ݜ����?�            pr@               
                     �?����˵�?O            �]@              	                 hލC@�\=lf�?.            �P@                                ���;@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        +            �N@                                   �?`�H�/��?!            �I@                                  �?؇���X�?            �A@                                 �*@�>����?             ;@                                 �B@ףp=
�?             4@       ������������������������       �                     1@                                  �'@�q�q�?             @        ������������������������       �                     �?                                   D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  �6@      �?              @                                ��m1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     0@               Q                     �?nS޸��?p             f@              P                 @�:x@�d�����?;            �W@              ?                    �?�5��
J�?9             W@              *                    �?R���Q�?'             N@                !                   �7@z�G�z�?             4@        ������������������������       �                     �?        "       )                 ��2>@�S����?             3@        #       (                    �?���Q��?             @       $       '                 ���<@      �?             @       %       &                   @@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        +       0                   �<@      �?             D@        ,       -                   �;@�q�q�?             @        ������������������������       �                     �?        .       /                 ��iB@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       >                    �?�L���?            �B@       2       =                   �>@�#-���?            �A@       3       4                 `fF:@R���Q�?             4@        ������������������������       �                     @        5       :                   @=@z�G�z�?	             .@       6       7                   `G@"pc�
�?             &@        ������������������������       �                     @        8       9                   @L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ;       <                   @K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             .@        ������������������������       �                      @        @       O                    �?     ��?             @@       A       B                 `fFJ@|��?���?             ;@        ������������������������       �                     @        C       N                 �U�X@\X��t�?             7@       D       E                    �?�����?             3@        ������������������������       �                     $@        F       M                 03�U@�q�q�?             "@       G       L                 `f�N@      �?              @       H       I                    7@      �?             @        ������������������������       �                     �?        J       K                    A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        R       U                    4@Ћ����?5            �T@        S       T                    &@�<ݚ�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        V       a                    �? �й���?1            @R@       W       `                    �?�O4R���?#            �J@       X       Y                   �)@p���?"             I@        ������������������������       �                     4@        Z       _                 �|�=@(;L]n�?             >@        [       \                 �|�<@��S�ۿ?
             .@       ������������������������       �                     $@        ]       ^                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     @        ������������������������       �                     4@        c       �                    @�����D�?�            `x@       d       e                    @tHN�?�             v@        ������������������������       �                     @        f       �                    �?*c̕6�?�            �u@        g       �                 �?�-@r�q��?>             X@       h       {                    �?l��
I��?2            @T@        i       z                 �� @     ��?             @@       j       k                    �?���N8�?             5@        ������������������������       �                     �?        l       y                 �|�=@z�G�z�?             4@       m       n                 ��y@����X�?	             ,@        ������������������������       �                      @        o       r                 ���@�q�q�?             (@        p       q                 �|�9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        s       t                   �<@�z�G��?             $@        ������������������������       �                     @        u       v                 �|Y=@և���X�?             @        ������������������������       �                     �?        w       x                   @@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        |       �                    �?`�(c�?            �H@        }       ~                 �|�9@�KM�]�?             3@        ������������������������       �                      @               �                    �?�t����?	             1@       �       �                  ��@      �?             0@        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     �?        �       �                  ��@��S�ۿ?             >@        ������������������������       �                     @        �       �                 ��(@���}<S�?             7@       �       �                 �|Y=@�����?             5@        ������������������������       �                     �?        �       �                 X��A@P���Q�?             4@       ������������������������       ��}�+r��?
             3@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?������?             .@       �       �                   �2@      �?              @        ������������������������       �                     �?        �       �                 ��$1@����X�?             @       �       �                    �?      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                    @      �?             @       �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �C@���S��?�            �o@       �       �                    �?|�5�L�?�            �k@        �       �                 @3�@X�Cc�?             E@        �       �                    �?      �?             (@       �       �                 pf�@�<ݚ�?             "@       ������������������������       �                     @        �       �                   �9@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 P�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?z�G�z�?             >@       �       �                 �|�;@����X�?             5@        �       �                    3@�C��2(�?             &@        �       �                 �y�+@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?      �?             $@       �       �                 �|�=@      �?             @        ������������������������       �                      @        �       �                    A@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 03�1@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        �       �                 �T)D@������?n            @f@       �       �                 �?�@t��ճC�?m             f@        �       �                    �?��
���?.            �R@       �       �                   �@��pBI�?,            @R@       �       �                 P�N@ �#�Ѵ�?            �E@       �       �                 ��@��Y��]�?            �D@       ������������������������       �                     <@        �       �                 �?$@$�q-�?             *@        �       �                 �|Y?@      �?              @       �       �                 �|Y8@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     >@        ������������������������       �                      @        �       �                 0SE @ܴD��??            @Y@        �       �                 ��) @z�G�z�?            �A@       �       �                    �?      �?             @@       �       �                 @3�@ 	��p�?             =@        �       �                   �A@r�q��?             @       ������������������������       �                     @        ������������������������       �      �?              @        �       �                   �3@�nkK�?             7@        �       �                   �1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     4@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    )@���7�?(            �P@        ������������������������       �                     �?        �       �                 `�X#@��ɉ�?'            @P@        �       �                    �?�FVQ&�?            �@@       �       �                 �|�=@`Jj��?             ?@       ������������������������       �                     6@        �       �                    ?@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @@        ������������������������       �                      @        ������������������������       �                     @@        �       �                    �?�X�<ݺ?             B@        ������������������������       �        
             1@        �       �                   �0@�KM�]�?             3@       �       �                 ��T?@��S�ۿ?             .@       ������������������������       �                     "@        �       �                    @r�q��?             @        �       �                 pf�C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������"N���I�?�c�~`l�?��j�F��?%�ʂ\��?              �?�}ylE��?W'u_�?��/���?W'u_�?g��1��?"=P9���?UUUUUU�?�������?              �?      �?                      �?�?�������?�$I�$I�?۶m۶m�?h/�����?�Kh/��?�������?�������?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?      �?      �?      �?      �?              �?      �?                      �?              �?G($��?�^o�?�?Cy�5��?y�5���?�,d!Y�?�Mozӛ�?333333�?333333�?�������?�������?              �?(������?^Cy�5�?�������?333333�?      �?      �?      �?      �?      �?                      �?              �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        }���g�?L�Ϻ��?�A�A�?_�_�?333333�?333333�?      �?        �������?�������?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?      �?              �?              �?      �?{	�%���?	�%����?      �?        ��Moz��?!Y�B�?^Cy�5�?Q^Cy��?              �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?              �?                      �?ԮD�J��?��+Q��?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?        ����Ǐ�?����?:�&oe�?�x+�R�?\���(\�?{�G�z�?      �?        �������?�?�������?�?      �?        �������?�������?      �?                      �?      �?              �?              �?        z�z��?z�z��?�2���?��5K�O�?              �?�֡�l�?Ȥx�L��?UUUUUU�?UUUUUU�?Lh/����?h/�����?      �?      �?�a�a�?��y��y�?              �?�������?�������?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?        ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?333333�?�������?      �?              �?              �?        ������?4և����?(�����?�k(���?              �?�?<<<<<<�?      �?      �?      �?                      �?      �?        �������?�?      �?        ӛ���7�?d!Y�B�?=��<���?�a�a�?              �?ffffff�?�������?�5��P�?(�����?      �?              �?        �?wwwwww�?      �?      �?      �?        �$I�$I�?�m۶m��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?      �?              �?      �?                      �?EQEQ�?]�u]�u�?�S�<%��?߰�k��?%I�$I��?�m۶m��?      �?      �?�q�q�?9��8���?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�m۶m��?�$I�$I�?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?              �?      �?              �?        ؽ�u�{�?B�P�"�?�E]t��?t�E]t�?&�X�%�?O贁N�?���Ǐ�?����?�/����?�}A_Ч?8��18�?������?      �?        �؉�؉�?;�;��?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?      �?      �?                      �?      �?              �?        �(0���?z��~�X�?�������?�������?      �?      �?������?�{a���?�������?UUUUUU�?      �?              �?      �?�Mozӛ�?d!Y�B�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�.�袋�?F]t�E�?              �??�?��? �����?>����?|���?���{��?�B!��?      �?        9��8���?�q�q�?              �?      �?              �?              �?                      �?      �?        ��8��8�?�q�q�?      �?        �k(���?(�����?�������?�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJڡWhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       j                     @�����?�           8�@               M                    �?&����j�?�            `t@                                  @���j��?�            �i@        ������������������������       �        	             0@               :                   �F@�ހ���?|            �g@                                  �?z91$UO�?\            �a@                                   �?�i�y�?)            �O@                                 �B@ �#�Ѵ�?            �E@       	                           9@P�Lt�<�?             C@        
                        ��*@@4և���?             ,@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     8@                                  �*@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@                                   $@H�z���?3             T@        ������������������������       �                      @               #                    �?����?1            �S@                                  �7@�q�q�?             ;@                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                ��";@�GN�z�?             6@        ������������������������       �                      @               "                    �?R���Q�?             4@              !                  Y>@�θ�?             *@                                 ���<@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        $       -                 ��$:@��x_F-�?"            �I@       %       *                   �@@��a�n`�?             ?@       &       )                    5@ ��WV�?             :@        '       (                    &@�8��8��?             (@        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �        
             ,@        +       ,                   @B@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        .       9                    �?��Q��?             4@       /       8                 ��yC@p�ݯ��?             3@       0       7                    D@���|���?             &@       1       4                 �|Y=@�z�G��?             $@        2       3                   @>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        5       6                   �>@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ;       B                    �?���X�K�?             �F@        <       =                    �?���!pc�?             &@        ������������������������       �                     �?        >       ?                     �?z�G�z�?             $@        ������������������������       �                     @        @       A                    L@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        C       L                   �R@��hJ,�?             A@       D       K                   �J@     ��?             @@       E       F                 `fF:@d}h���?             ,@        ������������������������       �                     @        G       J                 �T!@@      �?              @        H       I                   `G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                      @        N       [                    �?��6}��?H            �^@       O       R                    @`<)�+�?,            @S@        P       Q                 ��1V@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        S       T                    �?��pBI�?*            @R@        ������������������������       �                     9@        U       Z                    :@ �q�q�?             H@        V       Y                    �?؇���X�?
             ,@       W       X                   �E@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     A@        \       g                     �?�L�lRT�?            �F@        ]       f                    �?��Q��?             4@       ^       e                   �F@�����?             3@       _       `                 ��"@      �?
             0@        ������������������������       �                      @        a       b                  x#J@և���X�?	             ,@        ������������������������       �                     @        c       d                   �5@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        h       i                    (@H%u��?             9@        ������������������������       �                     @        ������������������������       �                     6@        k       �                    �?6��f�?�            x@       l       �                    �?z���=��?�            @s@        m       �                 ���1@�zv�X�?             F@       n       q                    3@�G�z�?             D@        o       p                 ��*@�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @        r       s                    5@� �	��?             9@        ������������������������       �                     �?        t       �                   @D@�q�q�?             8@       u       �                 �|�=@�û��|�?             7@       v       y                   �6@և���X�?             5@        w       x                 جJ"@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        z       �                 �?�@      �?             0@        {       |                 �|�<@      �?              @        ������������������������       �                     @        }       �                    �?      �?             @       ~                        �&�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                   �8@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �T)D@ ���]��?�            �p@       �       �                    �?��E���?�            `p@        �       �                   �6@x�����?            �C@        �       �                 ��y@�q�q�?             @        ������������������������       �                     �?        �       �                 �y.@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?<���D�?            �@@       �       �                 �|�;@��� ��?             ?@        �       �                   �8@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���@�>����?             ;@        ������������������������       �                     ,@        �       �                   @@8�Z$���?             *@        �       �                 �|�=@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�=�c��?�            �k@        �       �                 ��(@ �q�q�?             8@       �       �                 �|Y=@�X�<ݺ?             2@        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     @        �       �                   �7@�U6��?|            �h@        �       �                 @3�@�g�y��?)             O@       ������������������������       �                     @@        �       �                 0S5 @��S�ۿ?             >@        �       �                   �4@      �?              @       �       �                   �1@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     6@        �       �                 ��) @�6v��u�?S             a@       �       �                 @3�@�}�+r��?C            �\@       �       �                 �?�@���M�?4            @V@       �       �                 ���@������?.            �T@        ������������������������       �                     7@        �       �                 ���@ ,��-�?             �M@        ������������������������       �                      @        �       �                 �|Y=@���U�?            �L@        ������������������������       �                     9@        �       �                   @@@      �?             @@       �       �                   �@�KM�]�?             3@       �       �                 pf�@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     *@        �       �                   �?@����X�?             @        �       �                   �=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �A@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     9@        �       �                 ��y @��+7��?             7@        ������������������������       �                      @        �       �                    ?@��s����?             5@       �       �                   �:@�	j*D�?
             *@        ������������������������       �                     @        �       �                    �?      �?              @       �       �                    (@և���X�?             @       �       �                 ��)"@z�G�z�?             @        ������������������������       �                     �?        �       �                   �<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 �̌4@���|���?3            @S@        �       �                    �?     ��?             @@        �       �                 �|�:@և���X�?	             ,@       �       �                    �?؇���X�?             @       �       �                    &@      �?             @        ������������������������       �                      @        �       �                 83�0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    :@r�q��?             2@       ������������������������       �                     .@        ������������������������       �                     @        �       �                    @�����H�?            �F@        �       �                    �?�q�q�?	             (@        �       �                 @3;:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�z�G��?             $@       ������������������������       �                     @        �       �                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �B@Pa�	�?            �@@       ������������������������       �                     ;@        �       �                   �C@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub������������������?��܍��?!P�T��?p�W��(�?�?�������?      �?        ��Q�٨�?!&W�+�?�n��L�?��p��Y�?AA�?�������?�}A_Ч?�/����?(�����?���k(�?�$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?              �?�������?�������?      �?                      �?              �?�������?�������?              �?H�4H�4�?��-��-�?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?�袋.��?]t�E�?              �?333333�?333333�?ى�؉��?�؉�؉�?�$I�$I�?۶m۶m�?      �?                      �?      �?              �?        �������?�?�s�9��?�c�1Ƹ?O��N���?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        333333�?�������?UUUUUU�?UUUUUU�?      �?        �������?ffffff�?^Cy�5�?Cy�5��?F]t�E�?]t�E]�?333333�?ffffff�?      �?      �?      �?                      �?UUUUUU�?�������?              �?      �?              �?              �?              �?        l�l��?�'}�'}�?t�E]t�?F]t�E�?      �?        �������?�������?              �?�������?333333�?              �?      �?        KKKKKK�?�������?      �?      �?I�$I�$�?۶m۶m�?      �?              �?      �?      �?      �?      �?                      �?      �?              �?                      �?;ڼOq��?�!XG��?��O���?S{����?      �?      �?              �?      �?        ����?���Ǐ�?              �?UUUUUU�?�������?�$I�$I�?۶m۶m�?F]t�E�?/�袋.�?              �?      �?                      �?              �?�I��I��?l�l��?ffffff�?�������?^Cy�5�?Q^Cy��?      �?      �?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?              �?      �?        )\���(�?���Q��?              �?      �?        g�'�Y�?�cj`��?�cj`��?
qV~B��?�袋.��?��.���?�������?�������?�?�������?              �?      �?        )\���(�?�Q����?      �?        �������?�������?��,d!�?8��Moz�?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?      �?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?              �?      �?              �?        ���>��?>���>�?T���0�?�_�	)y�?��o��o�?�A�A�?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        |���?|���?�{����?�B!��?      �?      �?      �?                      �?�Kh/��?h/�����?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?333333�?�������?      �?              �?              �?        �������?xI@8�?�������?UUUUUU�?��8��8�?�q�q�?      �?      �?      �?                      �?      �?              �?        5q����?Zv<���?��{���?�B!��?      �?        �������?�?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?        c���s2�?�d�*al�?�5��P�?(�����?��^����?�E(B�?p>�cp�?������?      �?        [4���?'u_[�?              �?	�#����?p�}��?      �?              �?      �?�k(���?(�����?9��8���?�q�q�?      �?                      �?      �?              �?        �m۶m��?�$I�$I�?      �?      �?      �?                      �?�������?�������?      �?              �?      �?      �?        zӛ����?Y�B��?              �?z��y���?�a�a�?vb'vb'�?;�;��?      �?              �?      �?۶m۶m�?�$I�$I�?�������?�������?              �?      �?      �?      �?                      �?      �?              �?              �?                      �?]t�E]�?F]t�E�?      �?      �?۶m۶m�?�$I�$I�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?                      �?              �?�m۶m��?�$I�$I�?      �?                      �?UUUUUU�?�������?              �?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?ffffff�?333333�?      �?              �?      �?              �?      �?        |���?|���?      �?        �������?UUUUUU�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:d�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM'hjh))��}�(h,h/h0M'��h2h3h4hph<�h=Kub������       x                     @�4�O��?�           8�@                                   �?: �Z���?�            Pr@                                   �?H�̱���?Q            @_@        ������������������������       �                    �A@                                   6@�:�^���?:            �V@                                   L@���!pc�?             6@                                  �?�S����?             3@              	                 `f�)@      �?             0@        ������������������������       �                     @        
                           �?�C��2(�?             &@                                  ;@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                  �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �?г�wY;�?+             Q@        ������������������������       �                     ;@                                   �?������?            �D@                                  �C@؇���X�?             ,@                                   D@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ;@               =                    �?4և����?r             e@               <                   �H@�G�z��?             D@              ;                    �?��.k���?             A@              4                    �?�'�=z��?            �@@               1                    �?�\��N��?             3@       !       0                     �?և���X�?             ,@       "       +                   @@@      �?
             (@       #       &                  Y>@����X�?             @        $       %                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        '       (                 �M@z�G�z�?             @        ������������������������       �                     @        )       *                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ,       -                   �A@z�G�z�?             @        ������������������������       �                     @        .       /                 @�Cq@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        2       3                   �7@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        5       6                 ��G@և���X�?
             ,@        ������������������������       �                     @        7       8                   @H@z�G�z�?             $@        ������������������������       �                     @        9       :                 ���X@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        >       q                    �?     ��?T             `@       ?       b                     �?0y����?M            �]@        @       A                   �;@P̏����?&            �L@        ������������������������       �                      @        B       S                   �>@�rF���?$            �K@        C       R                    R@$��m��?             :@       D       Q                   �L@`�Q��?             9@       E       P                   �G@���Q��?             4@       F       G                 03:@�t����?
             1@        ������������������������       �                     @        H       I                 �|Y=@�eP*L��?             &@        ������������������������       �                      @        J       O                   @=@X�<ݚ�?             "@       K       L                 03k:@և���X�?             @        ������������������������       �                     �?        M       N                 `f�;@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        T       U                   @A@ܷ��?��?             =@        ������������������������       �        	             ,@        V       W                    �?z�G�z�?             .@        ������������������������       �                     @        X       Y                    D@      �?             (@        ������������������������       �                     �?        Z       _                    �?"pc�
�?             &@       [       ^                 �K@      �?              @        \       ]                  x#J@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        `       a                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        c       d                    �?�g�y��?'             O@        ������������������������       �                     �?        e       p                   �*@�]0��<�?&            �N@       f       i                    5@������?            �D@        g       h                   �2@r�q��?             @        ������������������������       �                     @        ������������������������       �      �?              @        j       k                   @D@��?^�k�?            �A@       ������������������������       �                     ;@        l       m                 `f�)@      �?              @        ������������������������       �                     @        n       o                   �F@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        r       w                 03c@X�<ݚ�?             "@       s       t                    �?����X�?             @        ������������������������       �                     �?        u       v                    1@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        y       �                  �#@v����?�             z@       z                          �0@.�ȓ�<�?�            �o@        {       |                    �?�eP*L��?             &@        ������������������������       �                     @        }       ~                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @@@J	9<���?�            `n@       �       �                    �?�46<�?~             i@        �       �                    �?\X��t�?"             G@       �       �                 P�*@v ��?             �E@        ������������������������       �                     �?        �       �                   �7@�G��l��?             E@        ������������������������       �                      @        �       �                 �|Y=@ҳ�wY;�?             A@        �       �                    �?���Q��?             @       �       �                   �<@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?8^s]e�?             =@        ������������������������       �                     @        �       �                 �|�=@�C��2(�?             6@       �       �                    �?�����?             5@        �       �                 ���@�����H�?             "@        ������������������������       �                     @        �       �                   @@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 ���@�8��8��?             (@        ������������������������       �                     �?        �       �                 ��(@�C��2(�?             &@       ������������������������       �ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �ٝ@؇���X�?\            @c@        ������������������������       �                     ;@        �       �                 �Yu@�h1�
U�?M            �_@        �       �                    �?�z�G��?             >@        �       �                    �?؇���X�?             @       �       �                 P��@z�G�z�?             @        ������������������������       �                      @        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        �       �                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��L@�LQ�1	�?             7@       ������������������������       �        	             1@        �       �                    =@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                 �?�@�*v��?;            @X@        ������������������������       �                     >@        �       �                 @3�@�'݊U�?*            �P@        �       �                    �?     ��?             0@       �       �                    �?      �?             ,@        �       �                   �9@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �?@      �?             $@       �       �                    :@X�<ݚ�?             "@       �       �                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�t����?"            �I@        �       �                 �|Y>@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?���H��?             E@       �       �                   �8@      �?             D@        �       �                   �3@�X�<ݺ?             2@       �       �                   �2@�����H�?             "@       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     "@        �       �                   �;@"pc�
�?             6@        ������������������������       �                     �?        �       �                 ��) @؇���X�?             5@       ������������������������       �        
             .@        �       �                 pf� @      �?             @        ������������������������       �                      @        �       �                 �|Y=@      �?             @        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 �?�@ �#�Ѵ�?            �E@       ������������������������       �                     <@        �       �                 @3�@�r����?             .@        ������������������������       �                      @        ������������������������       �        
             *@        �                           �?H�U?B�?[            �d@       �       �                    �?�;�vv��?/            @R@        �       �                    �?�c�Α�?             =@       �       �                    �?���B���?             :@        ������������������������       �                     @        �       �                    �?      �?
             4@       �       �                    �?�C��2(�?             &@        �       �                   �-@r�q��?             @       �       �                   �,@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ���.@X�<ݚ�?             "@        ������������������������       �                     @        �       �                 �|�;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @�X���?!             F@        �       �                    @����X�?	             ,@       �       �                    @      �?              @       �       �                    @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 `v�6@r�q��?             >@        �       �                   �/@���|���?
             &@       ������������������������       �                     @        ������������������������       �                     @        �       �                    @�}�+r��?             3@       ������������������������       �        
             *@        �       �                 ��T?@r�q��?             @        ������������������������       �                     @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?jJA��v�?,            �V@                                 7@���Q��?             $@        ������������������������       �                     @                              �0@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?                                 �?|��"J�?(            @T@                                @;@(N:!���?            �A@        	      
                   9@      �?              @       ������������������������       �                     @        ������������������������       �                      @                              �̬3@�>����?             ;@       ������������������������       �                     4@                                 �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @                                �*@��+7��?             G@        ������������������������       �                     @                                 �?R���Q�?             D@                              ��!>@      �?             @        ������������������������       �                     @        ������������������������       �                     �?              &                   @�8��8��?             B@                                �?ܷ��?��?             =@        ������������������������       �                     @                                 �?ȵHPS!�?             :@                                '@      �?             0@                              ��|2@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@               %                pf�C@ףp=
�?             $@       !      "                   @      �?             @        ������������������������       �                      @        #      $                ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M'KK��h2h3h4hVh<�h=Kub�������������X�>�?2�N����?L5���?A�Ye�	�?����Mb�?�ʡE���?              �?l�l��?}�'}�'�?t�E]t�?F]t�E�?^Cy�5�?(������?      �?      �?              �?F]t�E�?]t�E�?�q�q�?�q�q�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �?�?              �?������?p>�cp�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?%I�$I��?n۶m۶�?�������?�������?�?�������?|���?|��|�?y�5���?�5��P�?�$I�$I�?۶m۶m�?      �?      �?�m۶m��?�$I�$I�?      �?      �?      �?                      �?�������?�������?      �?              �?      �?      �?                      �?�������?�������?              �?      �?      �?      �?                      �?      �?        �������?333333�?              �?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?             ��?      �?�������?�5�5�??���#�?��Gp�?              �?yJ���?�־a��?�N��N��?vb'vb'�?��(\���?{�G�z�?333333�?�������?�������?�������?      �?        t�E]t�?]t�E�?      �?        �q�q�?r�q��?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?333333�?�������?      �?                      �?              �?      �?                      �?��=���?a���{�?      �?        �������?�������?      �?              �?      �?              �?/�袋.�?F]t�E�?      �?      �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?��{���?�B!��?      �?        \2�h��?;ڼOqɠ?p>�cp�?������?�������?UUUUUU�?      �?              �?      �?_�_��?�A�A�?      �?              �?      �?      �?        �������?�������?              �?      �?              �?        �q�q�?r�q��?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?              �?        B�eh��?|�4�/��?m6��f��?M&��d2�?]t�E�?t�E]t�?              �?�������?UUUUUU�?      �?                      �?��Ƭ4�?��L-�?H�z�G�?�z�G��?!Y�B�?��Moz��?G�w��?qG�w��?      �?        1�0��?��y��y�?              �?�������?�������?�������?333333�?      �?      �?      �?                      �?              �?|a���?	�=����?              �?]t�E�?F]t�E�?=��<���?�a�a�?�q�q�?�q�q�?      �?        �������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        ]t�E�?F]t�E�?�������?�������?      �?              �?              �?        ۶m۶m�?�$I�$I�?      �?        �N���t�?��b�X,�?ffffff�?333333�?�$I�$I�?۶m۶m�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?��Moz��?Y�B��?      �?              �?      �?      �?                      �?��Id��?�i�n�'�?      �?        ����?��[���?      �?      �?      �?      �?      �?      �?      �?                      �?      �?      �?�q�q�?r�q��?�$I�$I�?۶m۶m�?      �?                      �?              �?      �?              �?        <<<<<<�?�?�q�q�?�q�q�?      �?                      �?�0�0�?��y��y�?      �?      �?��8��8�?�q�q�?�q�q�?�q�q�?      �?              �?      �?      �?        /�袋.�?F]t�E�?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?      �?      �?      �?      �?                      �?      �?              �?        �/����?�}A_Ч?      �?        �������?�?              �?      �?        �D�JԮ�?�v%jW��?�8�?����Ǐ�?�{a���?5�rO#,�?ى�؉��?��؉���?              �?      �?      �?F]t�E�?]t�E�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�q�q�?r�q��?      �?        UUUUUU�?�������?      �?                      �?      �?        ]t�E�?�E]t��?�$I�$I�?�m۶m��?      �?      �?�������?�������?              �?      �?              �?                      �?�������?UUUUUU�?]t�E]�?F]t�E�?      �?                      �?�5��P�?(�����?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?        8�C8�C�?�����?�������?333333�?              �?�������?�������?      �?                      �?�E��ӭ�?�����H�?|�W|�W�?�A�A�?      �?      �?      �?                      �?�Kh/��?h/�����?      �?        �m۶m��?�$I�$I�?      �?                      �?zӛ����?Y�B��?              �?333333�?333333�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?��=���?a���{�?      �?        ��N��N�?�؉�؉�?      �?      �?333333�?�������?              �?      �?              �?        �������?�������?      �?      �?      �?              �?      �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�I]fhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM#hjh))��}�(h,h/h0M#��h2h3h4hph<�h=Kub������       �                 ��K.@�L*�<�?�           8�@              -                    �?����?�             x@               ,                   P,@�=���D�?9            �T@                                   @�w�"w��?5             S@                                `f�)@���}<S�?             7@        ������������������������       �                      @                                  �*@�r����?
             .@                                  B@"pc�
�?             &@       	                           �?ףp=
�?             $@       
                           :@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               '                    �?H(���o�?#            �J@                                  �?�q�q�?             H@                                ���@�KM�]�?             3@        ������������������������       �                     @                                   �?r�q��?	             (@        ������������������������       �                     �?                                   �?"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @                                ���@l��[B��?             =@        ������������������������       �                     @                                 `�X!@�q�q�?             8@                                 �9@؇���X�?             ,@       ������������������������       �                      @                                �|�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        !       &                   �8@z�G�z�?             $@        "       #                 �[$@���Q��?             @        ������������������������       �                      @        $       %                 ��&@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        (       +                    @���Q��?             @       )       *                    1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        .       �                    �?4�R�f�?�             s@       /       �                   @E@�1h�'��?�            `r@       0       1                 03�@$Z�?�            �p@        ������������������������       �                    �F@        2       �                   �D@�X�C�?�             l@       3       N                 �?$@L������?�            `k@        4       I                 ��@��d��?(            �O@       5       B                  ��@���5��?$            �L@       6       9                   �7@�L���?            �B@        7       8                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        :       A                 �Y�@�g�y��?             ?@        ;       <                 ���@$�q-�?	             *@        ������������������������       �                     @        =       >                 �|=@؇���X�?             @        ������������������������       �                     @        ?       @                 �|�=@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     2@        C       H                    �?z�G�z�?             4@       D       E                 �|Y=@���y4F�?
             3@        ������������������������       �                     �?        F       G                    �?r�q��?	             2@       ������������������������       �z�G�z�?             .@        ������������������������       �                     @        ������������������������       �                     �?        J       K                 �|Y8@      �?             @        ������������������������       �                      @        L       M                 �|Y?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        O       T                   �2@�:�^���?X            �c@        P       S                 pf� @����X�?             @        Q       R                    1@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        U       b                     @l������?S            �b@        V       W                   �(@������?            �B@        ������������������������       �                     &@        X       a                 ��,@8�Z$���?             :@       Y       ^                    @@"pc�
�?             6@       Z       ]                 �|�=@��S�ۿ?	             .@       [       \                 �|�<@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        _       `                   @B@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        c       r                 @3�@@4և���?@             \@        d       k                 �|Y=@�*/�8V�?            �G@        e       j                   �<@�㙢�c�?             7@       f       g                 �?�@�����?             5@       ������������������������       �        
             0@        h       i                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        l       m                    �? �q�q�?             8@        ������������������������       �                     @        n       o                    ?@�}�+r��?             3@       ������������������������       �                     .@        p       q                   �@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        s       t                   �<@P�2E��?#            @P@        ������������������������       �                     9@        u       �                    �?��(\���?             D@       v       w                 ��) @$�q-�?            �C@       ������������������������       �                     ;@        x       �                    ?@      �?	             (@       y       �                 �|�=@      �?             @       z       }                 �|Y=@���Q��?             @        {       |                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ~                        �̜&@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���%@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     9@        �       �                    �?�z�G��?             $@       �       �                    4@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �                         �R@H�5�E6�?�            Pt@       �       �                    B@ �qm���?�            �p@       �       �                   �@@�+�*��?x            �h@       �       �                    @�q�q�?S            �a@       �       �                    �?�b��-8�?H            �_@       �       �                    &@�nkK�?%            @Q@        �       �                    �?�����H�?             2@       �       �                    �?"pc�
�?             &@       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��.@���J��?            �I@        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �H@        �       �                    �?F�����?#            �L@       �       �                    �?�û��|�?              G@       �       �                 ��$:@h+�v:�?             A@       �       �                 �|=@�t����?             1@        ������������������������       �                     @        �       �                  �v6@z�G�z�?             $@       ������������������������       �                     @        �       �                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?ҳ�wY;�?             1@       �       �                    <@������?
             .@        ������������������������       �                     @        �       �                 `f&;@���Q��?             $@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                 �|�?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �<@���Q��?             @        ������������������������       �                     �?        �       �                 �|Y=@      �?             @        ������������������������       �                     �?        �       �                   �>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?             (@        ������������������������       �                     @        �       �                 039@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?���!pc�?             &@        ������������������������       �                     @        �       �                    +@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�r����?             .@        ������������������������       �                     @        �       �                 �|Y?@"pc�
�?             &@       �       �                    @ףp=
�?             $@       �       �                 ��T?@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                     @h�����?%             L@       �       �                    �?     ��?             @@       �       �                    �?�G�z��?             4@       �       �                 03�J@�q�q�?	             (@       ������������������������       �                     @        �       �                     �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   PP@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �D C@r�q��?	             (@        �       �                    0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?ףp=
�?             $@       ������������������������       �                      @        �       �                     �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?r�q��?             8@        �       �                    ;@z�G�z�?             @        ������������������������       �                     @        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        �       �                    �?^H���+�?/            �R@        �       �                    @�GN�z�?             6@       �       �                    �?��s����?             5@        �       �                   �H@      �?             (@        ������������������������       �                     @        �       �                     �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @�����H�?             "@       ������������������������       �                     @        �       �                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?D>�Q�?"             J@        �       �                    �?z�G�z�?             $@       �       �                 pV�F@���Q��?             @       �       �                 p�i@@      �?             @       �       �                 ��Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                   �?r�q��?             E@                                R@�������?             >@                                �?V�a�� �?             =@             
                  �J@���N8�?             5@             	                �T!@@�eP*L��?             &@                               �G@      �?              @                                 G@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@                              �K@      �?              @                               x#J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@                                 �?�{��?��?&             K@                              "�b@��?^�k�?            �A@       ������������������������       �                     7@                                 �?�8��8��?             (@        ������������������������       �                     @                              Ъ�c@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @              "                   �?�\��N��?             3@             !                �̾w@     ��?             0@                              03c@�q�q�?
             (@                               �D@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M#KK��h2h3h4hVh<�h=Kub������������KY� ��?iM���{�?���H	�?�T�/���?�+Q��?w%jW�v�?��k(��?���k(�?d!Y�B�?ӛ���7�?              �?�?�������?F]t�E�?/�袋.�?�������?�������?      �?      �?      �?                      �?              �?      �?                      �?e�Cj���?M0��>��?UUUUUU�?UUUUUU�?(�����?�k(���?              �?UUUUUU�?�������?              �?F]t�E�?/�袋.�?              �?      �?        GX�i���?���=��?              �?�������?�������?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?333333�?�������?      �?      �?              �?      �?                      �?      �?        (������?����k�?K���+�?�E�_���?ɡ.K5��?��U��?      �?        �$I�$I�?n۶m۶�?�Ǐ?~�?����?��뺮��?EQEQ�?�}��?��Gp�?}���g�?L�Ϻ��?UUUUUU�?UUUUUU�?              �?      �?        ��{���?�B!��?�؉�؉�?;�;��?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        �������?�������?6��P^C�?(������?              �?�������?UUUUUU�?�������?�������?      �?              �?              �?      �?      �?              �?      �?              �?      �?        � � �?�o��o��?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        +�3�=l�?��c.��?��g�`��?к����?      �?        ;�;��?;�;��?/�袋.�?F]t�E�?�������?�?۶m۶m�?�$I�$I�?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?              �?        n۶m۶�?�$I�$I�?r1����?m�w6�;�?�7��Mo�?d!Y�B�?=��<���?�a�a�?      �?        333333�?�������?      �?                      �?              �?�������?UUUUUU�?      �?        �5��P�?(�����?      �?              �?      �?              �?      �?        _�^��?z�z��?      �?        �������?333333�?�؉�؉�?;�;��?      �?              �?      �?      �?      �?333333�?�������?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?        ffffff�?333333�?�$I�$I�?۶m۶m�?              �?      �?              �?        �t|��?�������?	��3���?��f,�?���W�?	��wT�?UUUUUU�?UUUUUU�?QEQE�?�u]�u]�?d!Y�B�?�Mozӛ�?�q�q�?�q�q�?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�?______�?      �?      �?              �?      �?                      �?u�YLg�?�YLg1�?8��Moz�?��,d!�?�������?xxxxxx�?<<<<<<�?�?      �?        �������?�������?      �?              �?      �?      �?                      �?�������?�������?�?wwwwww�?              �?�������?333333�?�������?�������?              �?      �?      �?      �?                      �?333333�?�������?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?              �?9��8���?�q�q�?      �?                      �?t�E]t�?F]t�E�?              �?333333�?�������?              �?      �?        �������?�?      �?        /�袋.�?F]t�E�?�������?�������?�������?�������?      �?                      �?      �?                      �?n۶m۶�?%I�$I��?      �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?              �?      �?              �?      �?        UUUUUU�?�������?      �?      �?              �?      �?        �������?�������?              �?      �?      �?              �?      �?        �������?UUUUUU�?�������?�������?              �?      �?      �?      �?                      �?      �?        L�Ϻ��?�g�`�|�?]t�E�?�袋.��?�a�a�?z��y���?      �?      �?              �?      �?      �?      �?                      �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        b'vb'v�?vb'vb'�?�������?�������?333333�?�������?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?        �������?UUUUUU�?�������?�������?��{a�?a���{�?�a�a�?��y��y�?t�E]t�?]t�E�?      �?      �?      �?      �?      �?      �?      �?                      �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        /�����?���^B{�?�A�A�?_�_��?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?      �?                      �?y�5���?�5��P�?      �?      �?�������?�������?      �?      �?              �?      �?              �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�޵#hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM;hjh))��}�(h,h/h0M;��h2h3h4hph<�h=Kub������       
                 x#J@"��p�?�           8�@              ]                 `f�$@������?r           ��@                                   �?�O~�B�?�            �p@                                   �?�q�q�?/            �S@               
                 ���@�������?             A@                                03S@@4և���?	             ,@        ������������������������       �                      @               	                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@                                  �5@���Q��?             4@        ������������������������       �                     @                                �|Y=@z�G�z�?             .@                                  @@      �?             @       ������������������������       �                      @        ������������������������       �                      @                                �|�=@�C��2(�?             &@                               p&�@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?�zv�X�?             F@                                   �?��s����?             5@                               ���@�X�<ݺ?
             2@        ������������������������       �                     �?        ������������������������       �        	             1@        ������������������������       �                     @        ������������������������       �                     7@               \                    �?���[�A�?|             h@              %                    �?����{�?{            �g@               $                    �?      �?             8@               !                   �@և���X�?             5@        ������������������������       �                      @        "       #                    4@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @        &       S                 ���"@�-�����?n            �d@       '       (                     @@݈g>h�?e             c@        ������������������������       �                     "@        )       N                    �?�C����?_            �a@       *       5                 P�N@     �?W             `@        +       ,                 ���@h㱪��?!            �K@        ������������������������       �                     7@        -       .                 ���@      �?             @@        ������������������������       �                     �?        /       0                 ��@�g�y��?             ?@        ������������������������       �        	             ,@        1       2                 �|�<@�IєX�?             1@       ������������������������       �                     &@        3       4                 �|Y>@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        6       9                 �Yu@0�й���?6            @R@        7       8                    >@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        :       C                    ?@t�e�í�?3            �P@       ;       B                   �3@ ��WV�?'             J@        <       =                 �?�@�<ݚ�?             "@        ������������������������       �                     @        >       ?                   �1@���Q��?             @        ������������������������       �                      @        @       A                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                    �E@        D       I                   �@@z�G�z�?             .@        E       F                 �?�@�q�q�?             @        ������������������������       �                     �?        G       H                 ��I @���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        J       K                   @C@�����H�?             "@        ������������������������       �                     @        L       M                 @3�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        O       P                 P�@z�G�z�?             .@       ������������������������       �                     "@        Q       R                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        T       U                   �<@���Q��?	             .@       ������������������������       �                     @        V       [                   �?@      �?              @       W       Z                 �|�=@؇���X�?             @       X       Y                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ^                       `f�C@��}*$&�?�            Pt@       _       l                    @Tt�ó��?�            `r@        `       a                     @��� ��?             ?@        ������������������������       �                     *@        b       c                    @�<ݚ�?             2@       ������������������������       �                     "@        d       g                    �?X�<ݚ�?             "@        e       f                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        h       i                    �?      �?             @        ������������������������       �                     �?        j       k                    @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        m       �                   �A@�:)<Q��?�            pp@       n       �                 �B,@�����?l            �e@        o       x                    �?�������?#             N@        p       q                    �?h�����?             <@        ������������������������       �                     "@        r       s                 ��y)@�}�+r��?
             3@        ������������������������       �                     "@        t       w                    �?ףp=
�?             $@       u       v                    :@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        y       z                    .@      �?             @@        ������������������������       �                      @        {       �                    �?��S�ۿ?             >@       |       }                 `fF)@�>����?             ;@        ������������������������       �                     $@        ~                           @@�t����?	             1@       ������������������������       �                     .@        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��K.@�Cc}h,�?I             \@        �       �                    �?�r����?
             .@       �       �                   �0@�C��2(�?             &@        �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 `f�,@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    '@�d�~V��??            @X@        �       �                     @r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        �       �                     @Zz�����?8            @U@       �       �                   �<@#z�i��?            �D@        �       �                    �?@�0�!��?             1@        ������������������������       �                     @        �       �                    �?d}h���?             ,@       �       �                    �?ףp=
�?             $@        �       �                   @<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?             @       �       �                   �7@�q�q�?             @        ������������������������       �                     �?        �       �                   �:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     �?r�q��?             8@       �       �                 �|�?@��
ц��?	             *@       �       �                 �|Y=@���|���?             &@        ������������������������       �                      @        �       �                    �?X�<ݚ�?             "@        �       �                 ��2>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   `@@      �?             @       �       �                 `f�<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �D`A@���|���?             &@       �       �                   @=@�z�G��?             $@       �       �                   �?@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?���|���?             F@        �       �                    �?�<ݚ�?             2@       �       �                    �?     ��?	             0@        ������������������������       �                     @        �       �                 03�3@�z�G��?             $@       �       �                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?$�q-�?             :@        �       �                 @34@z�G�z�?             $@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             0@        �       �                    �?�����?5            �V@       �       �                    �?:���W�?#            �M@        �       �                    �?�S����?
             3@       �       �                    D@      �?             0@        ������������������������       �                     �?        �       �                   �'@��S�ۿ?             .@        �       �                   �J@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                     �?�q�q�?             @        ������������������������       �                     �?        �       �                 03�5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             D@        �       �                 p�i@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�L���?            �B@       �       �                     �?l��\��?             A@        �       �                  )?@�r����?
             .@       �       �                    R@      �?              @       �       �                   �J@؇���X�?             @        �       �                   �H@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @�}�+r��?             3@       �       �                   �*@�IєX�?             1@       �       �                 `f�)@      �?              @        ������������������������       �                      @        �       �                    G@r�q��?             @        �       �                   �C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        �       �                     @     ��?             @@        �       �                    �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��T?@�����?             5@       ������������������������       �        
             2@        �                        ��p@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 I@��� ��?             ?@                                @ܷ��?��?             =@                               �8@r�q��?             2@        ������������������������       �                     @        ������������������������       �        	             .@        ������������������������       �                     &@              	                 �>I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              p�1N@��VT4�?I            �\@                              `fK@      �?             8@                                 �?      �?              @                                7@����X�?             @        ������������������������       �                     �?                                 �?r�q��?             @        ������������������������       �                      @                              `�iJ@      �?             @        ������������������������       �                     �?                                 @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                   @      �?	             0@       ������������������������       �                     &@                              �|�;@z�G�z�?             @        ������������������������       �                     @                              �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              :                   @�	j*D�?9            �V@              !                ��UO@ι�~��?5            �U@        ������������������������       �                     @        "      9                  �L@���Fi�?3            �T@       #      2                   �?���B���?0            �S@       $      )                �|Y<@��|�5��?            �G@        %      &                   �?���Q��?	             .@        ������������������������       �                     @        '      (                 �}S@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        *      +                  �D@     ��?             @@        ������������������������       �        	             .@        ,      -                   �?�t����?	             1@        ������������������������       �                      @        .      /                   G@X�<ݚ�?             "@        ������������������������       �                     �?        0      1                @�pX@      �?              @        ������������������������       �                     @        ������������������������       �                     @        3      8                   �?��� ��?             ?@       4      5                   �?���y4F�?             3@       ������������������������       �        	             ,@        6      7                  �G@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M;KK��h2h3h4hVh<�h=Kub������������J54v��?l�����?�?��8��?܀�����?�ݛ�D�?���)��?UUUUUU�?UUUUUU�?�������?�������?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?              �?�������?�������?      �?      �?      �?                      �?]t�E�?F]t�E�?�������?UUUUUU�?�������?�������?      �?              �?        ��.���?�袋.��?�a�a�?z��y���?�q�q�?��8��8�?      �?                      �?      �?              �?        %�T�/��?ko��@��?��U@0$�?,��>o�?      �?      �?�$I�$I�?۶m۶m�?              �?�؉�؉�?;�;��?              �?      �?              �?        u,e�*�?\��l���?�P^Cy�?Cy�5��?      �?        T�ik���?_���?     @�?      �?־a���?��)A��?      �?              �?      �?              �?��{���?�B!��?      �?        �?�?      �?        �������?UUUUUU�?      �?      �?      �?        ����?����Ǐ�?UUUUUU�?UUUUUU�?      �?                      �?�1����?�rv��?O��N���?;�;��?9��8���?�q�q�?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?      �?      �?        �q�q�?�q�q�?      �?              �?      �?              �?      �?        �������?�������?      �?              �?      �?              �?      �?        333333�?�������?      �?              �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?&�5����?�ߔ���?h�����?/�����?�B!��?�{����?              �?�q�q�?9��8���?              �?�q�q�?r�q��?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?        �������?333333�?              �?      �?        ���m9�?ɾ�$��?_��}�?A_���?�������?�������?�$I�$I�?�m۶m��?              �?(�����?�5��P�?              �?�������?�������?�$I�$I�?۶m۶m�?      �?                      �?              �?      �?      �?              �?�������?�?�Kh/��?h/�����?      �?        <<<<<<�?�?      �?                      �?      �?        %I�$I��?�m۶m��?�������?�?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?              �?      �?      �?              �?      �?      �?                      �?�i�n�'�?�,O"Ӱ�?�������?UUUUUU�?              �?      �?        �������?000000�?ە�]���?�+Q��?�������?ZZZZZZ�?              �?۶m۶m�?I�$I�$�?�������?�������?      �?      �?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?�;�;�?�؉�؉�?]t�E]�?F]t�E�?      �?        r�q��?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?      �?                      �?      �?                      �?F]t�E�?]t�E]�?333333�?ffffff�?      �?      �?              �?333333�?�������?              �?      �?                      �?      �?        ]t�E]�?F]t�E�?�q�q�?9��8���?      �?      �?              �?333333�?ffffff�?�$I�$I�?�m۶m��?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �؉�؉�?;�;��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        h�h��?�/��/��?_[4��?A�Iݗ��?^Cy�5�?(������?      �?      �?      �?        �?�������?�������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?        }���g�?L�Ϻ��?------�?�������?�������?�?      �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �5��P�?(�����?�?�?      �?      �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?              �?              �?      �?]t�E]�?F]t�E�?              �?      �?        =��<���?�a�a�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �{����?�B!��?��=���?a���{�?�������?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?m5x�@�?vI�ø_�?      �?      �?      �?      �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?�������?�������?              �?      �?      �?      �?                      �?;�;��?vb'vb'�?G�w��?�w�q�?      �?        ��FS���?�C.+J�?ى�؉��?��؉���?x6�;��?br1���?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?�������?�������?              �?r�q��?�q�q�?      �?              �?      �?              �?      �?        �B!��?�{����?(������?6��P^C�?              �?�������?�������?      �?                      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�G�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       .                   �1@�t����?�           8�@                                    @�X���?@             \@               
                     �?�#-���?            �A@                                   �?�z�G��?             $@        ������������������������       �                     @                                ��f`@���Q��?             @        ������������������������       �                     �?               	                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     9@               !                    @�eP*L��?,            @S@                                  �?(���@��?            �G@                                 �0@f.i��n�?            �F@                               03�-@�MI8d�?            �B@                                  /@�>����?             ;@       ������������������������       �        	             4@                                   �?����X�?             @        ������������������������       �                     @                                pf�@      �?             @        ������������������������       �                     �?                                �̌!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   #@���Q��?             $@                                  �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        "       -                    @ףp=
�?             >@       #       $                    �?�LQ�1	�?             7@        ������������������������       �                     (@        %       &                    @���!pc�?             &@        ������������������������       �                     @        '       ,                    �?      �?              @       (       )                 ���3@����X�?             @        ������������������������       �                     �?        *       +                    @r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        /       p                    �?���\˾�?           ��@        0       =                     @8�f�ȭ�?�            `h@       1       <                    �? ;=֦��?L            �^@       2       3                   �H@ �q�q�?-             R@       ������������������������       �        %             M@        4       ;                 ,w�U@d}h���?             ,@       5       :                   �L@�q�q�?             "@       6       9                    L@      �?              @       7       8                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     I@        >       Q                    �?�6����?4            @R@        ?       P                    �?      �?             @@       @       G                    �?���Q��?             4@        A       B                   �7@      �?             @        ������������������������       �                      @        C       D                 X�x&@      �?             @        ������������������������       �                     �?        E       F                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        H       O                 03@X�Cc�?
             ,@       I       J                 �|�9@      �?             $@        ������������������������       �                     �?        K       N                    �?X�<ݚ�?             "@       L       M                  ��@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        R       o                   �C@��]�T��?             �D@       S       b                    �?�q�q�?             B@       T       _                   �;@j���� �?             1@       U       ^                    �?�	j*D�?             *@       V       [                 pf� @���|���?
             &@       W       Z                   �3@؇���X�?             @        X       Y                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        \       ]                  �#@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        `       a                 pf�$@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        c       n                    @�d�����?             3@       d       e                 �|Y=@�<ݚ�?             2@        ������������������������       �                     "@        f       m                   �>@X�<ݚ�?             "@       g       l                     @      �?              @       h       k                 �|�=@      �?             @       i       j                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        q       �                     �?�Mc��?�            @y@        r                           �?T��o��?;            @W@        s       |                    �?���!pc�?            �@@       t       {                 �̾w@�㙢�c�?             7@       u       z                    �?�����?             5@       v       y                 �|Y<@�r����?
             .@        w       x                  �}S@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                      @        }       ~                 �UcV@      �?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�0u��A�?$             N@       �       �                   �<@>n�T��?#             M@        �       �                    �?8�Z$���?             *@       ������������������������       �                     $@        �       �                    7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �G@������?            �F@       �       �                 ��<:@6YE�t�?            �@@        ������������������������       �                     @        �       �                 �T!@@�>4և��?             <@        �       �                   �C@�q�q�?             "@       �       �                 `f�<@���Q��?             @       �       �                 �|�?@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y>@�KM�]�?             3@        ������������������������       �                     "@        �       �                  x#J@z�G�z�?             $@        ������������������������       �                     @        �       �                    A@�q�q�?             @        ������������������������       �                     �?        �       �                 `�iJ@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             (@       �       �                   @L@X�<ݚ�?             "@        ������������������������       �                     @        �       �                 `fF<@r�q��?             @       ������������������������       �                     @        �       �                  )?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?0��O�?�            ps@        �       �                   �6@�3Ea�$�?             G@        �       �                    �?r�q��?             @       �       �                    5@z�G�z�?             @       �       �                 �{@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?ףp=
�?             D@       �       �                 �|Y=@��� ��?             ?@        �       �                   �<@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�=@ �q�q�?             8@       �       �                 ���@�X�<ݺ?
             2@        ������������������������       �                     @        �       �                   @@�8��8��?             (@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �                          �?��ckݭ�?�            �p@       �       �                    �?���Lͩ�?�             l@        �       �                     @P���Q�?             4@        ������������������������       �                     �?        �       �                 X��A@�}�+r��?             3@       �       �                 �Y�@��S�ۿ?
             .@        ������������������������       �                     @        ������������������������       ��8��8��?             (@        ������������������������       �                     @        �                          �?������?�            �i@       �       �                   �<@����#��?~             i@        �       �                 ���@���N8�?6             U@        �       �                 ���@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                     @�g<a�?2            @S@        �       �                    &@��S�ۿ?
             .@        �       �                   �5@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �3@0�z��?�?(             O@        �       �                 �?�@$�q-�?	             *@       ������������������������       �                      @        �       �                 0S5 @z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                    �H@        �                        0��D@�����8�?H            @]@       �       �                     @d�X^_�?G            �\@        �       �                   @F@������?            �D@       �       �                 `fF)@\-��p�?             =@        ������������������������       �                     *@        �       �                   �3@      �?             0@       �       �                 �|�=@���|���?             &@        ������������������������       �                      @        �       �                   @D@�<ݚ�?             "@       �       �                    @@      �?              @        ������������������������       �                     @        �       �                   @B@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                   @@@$G$n��?0            �R@       �       �                 �|Y>@��P���?            �D@       �       �                 �|Y=@ܷ��?��?             =@        �       �                 ���"@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                  sW@�8��8��?             8@        �       �                 ��,@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     .@        �       �                   �?@      �?             (@        ������������������������       �                     �?        �       �                   �@�eP*L��?             &@        ������������������������       �                     @        �       �                 �?�@      �?              @        ������������������������       �                     �?        �       �                 ��I @����X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                 @3�@Pa�	�?            �@@       �       �                 �?�@      �?             0@       ������������������������       �                     ,@        ������������������������       �      �?              @        ������������������������       �                     1@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     D@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������G�+J>�?r%�k���?n۶m۶�?I�$I�$�?_�_�?�A�A�?333333�?ffffff�?              �?333333�?�������?              �?      �?      �?      �?                      �?              �?t�E]t�?]t�E�?R�٨�l�?W�+���?�>�>��?�`�`�?L�Ϻ��?��L���?h/�����?�Kh/��?              �?�$I�$I�?�m۶m��?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?      �?      �?      �?                      �?      �?              �?              �?      �?              �?      �?        �������?�������?��Moz��?Y�B��?      �?        F]t�E�?t�E]t�?      �?              �?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?              �?      �?                      �?      �?        ��@?�?�:z�~��?��I��I�?ڞ�ٞ��?XG��).�?�%C��6�?UUUUUU�?�������?              �?۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?      �?      �?�$I�$I�?�m۶m��?      �?                      �?      �?                      �?              �?              �?�ܹs���?�#F��?      �?      �?�������?333333�?      �?      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?%I�$I��?      �?      �?              �?r�q��?�q�q�?�������?�������?      �?                      �?      �?                      �?              �?KԮD�J�?jW�v%j�?�������?�������?ZZZZZZ�?�������?;�;��?vb'vb'�?F]t�E�?]t�E]�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?Cy�5��?y�5���?9��8���?�q�q�?      �?        r�q��?�q�q�?      �?      �?      �?      �?      �?      �?              �?      �?              �?              �?                      �?              �?      �?        5r���?+�7����?���O?��?X`��?F]t�E�?t�E]t�?�7��Mo�?d!Y�B�?=��<���?�a�a�?�������?�?      �?      �?              �?      �?              �?              �?                      �?      �?      �?              �?      �?        �������?�������?,�4�rO�?��{a�?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?                      �?wwwwww�?�?'�l��&�?e�M6�d�?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?�������?333333�?      �?      �?      �?                      �?              �?      �?        �k(���?(�����?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?        �������?�������?r�q��?�q�q�?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        ˿!a���?���̱�?����7��?��,d!�?UUUUUU�?�������?�������?�������?      �?      �?      �?                      �?              �?              �?�������?�������?�{����?�B!��?�$I�$I�?۶m۶m�?      �?                      �?�������?UUUUUU�?��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?              �?              �?        ZK���v�?1��:kI�?�6�i�?�K~��?ffffff�?�������?      �?        �5��P�?(�����?�������?�?      �?        UUUUUU�?UUUUUU�?      �?        �|����?������?���(���?�C��x�?��y��y�?�a�a�?�m۶m��?�$I�$I�?      �?                      �?���8+�?�cj`?�������?�?�������?�������?      �?      �?      �?              �?        |���{�?�B!��?�؉�؉�?;�;��?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?        �������?���?�s���?�aܯK*�?�|����?������?a����?�{a���?      �?              �?      �?]t�E]�?F]t�E�?              �?9��8���?�q�q�?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        к����?���L�?������?�����?��=���?a���{�?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?9��8���?�q�q�?      �?                      �?      �?              �?      �?              �?t�E]t�?]t�E�?              �?      �?      �?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?        |���?|���?      �?      �?      �?              �?      �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���JhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM#hjh))��}�(h,h/h0M#��h2h3h4hph<�h=Kub������       �                     @���;+"�?�           8�@               m                    �? Q�TG�?�            v@              F                     �?�Z����?�             q@               3                 ��9L@~�hP��?N            �b@              
                    �?      �?.            �T@               	                 03�=@�C��2(�?
             6@                                ���;@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@                                   �?��Q��?$             N@                                �|�;@������?	             .@        ������������������������       �                     �?                                p�i@@d}h���?             ,@                               ���<@�q�q�?             "@        ������������������������       �                     @                                  �H@      �?             @                               X�lA@���Q��?             @                               ��2>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               2                   @L@F�����?            �F@              -                    �?H�z�G�?             D@              ,                   �G@�ʻ����?             A@              +                 ��yC@J�8���?             =@                               ��I*@      �?             4@        ������������������������       �                     @                                 03k:@j���� �?             1@        ������������������������       �                      @        !       "                 �|�<@��S���?
             .@        ������������������������       �                     @        #       *                   �C@�z�G��?             $@       $       )                 �|�?@      �?             @       %       &                 `f�<@���Q��?             @        ������������������������       �                      @        '       (                   `@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        .       /                   �C@�q�q�?             @        ������������������������       �                     @        0       1                    G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        4       A                   �D@��2(&�?             �P@       5       @                    �?l�b�G��?            �L@       6       ?                 �|�=@�����H�?             B@       7       8                    �?z�G�z�?             4@       ������������������������       �                     *@        9       <                    �?և���X�?             @        :       ;                 �|Y<@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        =       >                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �        
             5@        B       E                 `f^@X�<ݚ�?             "@       C       D                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        G       H                    @b����?N            �_@        ������������������������       �                     $@        I       V                    �?����"�?J             ]@        J       O                    �?�C��2(�?             F@       K       N                   �:@�>����?             ;@        L       M                   �7@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     4@        P       U                   �E@�t����?             1@       Q       T                   �6@      �?             0@        R       S                 ��m1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                     �?        W       l                    ,@�X�<ݺ?/             R@       X       Y                    �?�8��8��?             H@        ������������������������       �                     �?        Z       _                 `f�)@dP-���?            �G@        [       ^                    &@ �q�q�?             8@       \       ]                    5@P���Q�?             4@        ������������������������       ��q�q�?             @        ������������������������       �        
             1@        ������������������������       �                     @        `       a                 �|�<@�LQ�1	�?             7@        ������������������������       �                     @        b       c                 �|�=@     ��?
             0@        ������������������������       �                     �?        d       e                    @@�r����?	             .@        ������������������������       �                     @        f       g                   �A@r�q��?             (@        ������������������������       �      �?              @        h       i                   @D@ףp=
�?             $@        ������������������������       �                     @        j       k                   �F@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     8@        n       s                    �?�6i����?.            �S@        o       p                   �7@�G��l��?             5@        ������������������������       �                     "@        q       r                    �?r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        t       }                    Q@\-��p�?"             M@       u       v                   �A@������?            �D@       ������������������������       �                     @@        w       x                    �?�<ݚ�?             "@        ������������������������       �                     �?        y       |                     @      �?              @       z       {                    F@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ~       �                   @K@ҳ�wY;�?	             1@              �                 Ъ�c@8�Z$���?             *@        �       �                    �?      �?             @       �       �                    3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                    �?�K�J���?�            `v@        �       �                    �?��S���?B            @Z@       �       �                 03�0@&:~�Q�?0             S@       �       �                   �C@�c�Α�?%             M@       �       �                   �3@x��}�?$            �K@        �       �                 P��+@�IєX�?             1@       ������������������������       �        	             .@        �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y=@�����?             C@        �       �                   �;@�G��l��?             5@       �       �                 ��@X�<ݚ�?	             2@        ������������������������       �                     @        �       �                 ��&@���!pc�?             &@       �       �                   �9@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�IєX�?             1@       ������������������������       �                     &@        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�7@b�2�tk�?             2@        �       �                    �?"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                 �|Y>@����X�?             @       �       �                    @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?>���Rp�?             =@        �       �                    @      �?             @       �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?z�G�z�?             9@        ������������������������       �                     @        �       �                   �0@�GN�z�?             6@        ������������������������       �                     "@        �       �                 ��p@@�n_Y�K�?	             *@        �       �                    @r�q��?             @        ������������������������       �                     @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����sV�?�            �o@        �       �                 �|Y=@�E��ӭ�?             B@        �       �                 �&�)@�eP*L��?             &@       �       �                    ;@      �?              @       �       �                    0@���Q��?             @        ������������������������       �                      @        �       �                    5@�q�q�?             @        ������������������������       �                     �?        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�J�4�?             9@       �       �                 ���@���7�?             6@        ������������������������       �                     &@        �       �                   @@�C��2(�?             &@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        �                          @��� ��?�             k@       �       �                    �?      �?~             i@        �       �                    �? 7���B�?             ;@       �       �                    �? ��WV�?             :@       �       �                 �|Y;@�IєX�?             1@        ������������������������       �                     �?        �       �                 ���@      �?             0@        ������������������������       �                     @        �       �                 ��(@$�q-�?	             *@       ������������������������       ��C��2(�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        �                          �?E�Vl��?m            �e@       �       �                   �0@ףp=��?d             d@        �       �                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �9@P5�޷�?b            �c@        �       �                 ���@h㱪��?$            �K@        �       �                    7@�����H�?             "@       ������������������������       �                     @        �       �                   �8@z�G�z�?             @       �       �                 �&b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��<b�ƥ?             G@       ������������������������       �                     D@        �       �                 ��Y@r�q��?             @        ������������������������       �                     @        �       �                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �                       �T)D@��hJ,�?>            �Y@       �                          �?<���D�?=            �X@       �       �                   �;@H�g�}N�?9            �V@        �       �                   �:@�z�G��?             $@       ������������������������       �                     @        �       �                 �� @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �                         �C@�����H�?4            @T@       �                         @C@      �?-             R@       �                         @@@���Ls�?*            @P@       �                       �Yu@ȵHPS!�?"             J@        �                         �?@���|���?             &@                              ��@�z�G��?             $@        ������������������������       �                      @                              �&B@      �?              @                             �|Y>@և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                 ?@������?            �D@       	      
                ���"@P�Lt�<�?             C@       ������������������������       �                     @@                                 (@r�q��?             @                              �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     *@                              ��	0@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @                                 4@�n_Y�K�?	             *@                                  @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 �?@�0�!��?
             1@       ������������������������       �                     $@              "                   @և���X�?             @              !                   @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0M#KK��h2h3h4hVh<�h=Kub������������D�#{��?x��	��?MV)'
2�?�Tk��f�?�J���?��s2}��?�Y7�"��?S�n0�?      �?      �?F]t�E�?]t�E�?�������?�������?              �?      �?                      �?�������?ffffff�?wwwwww�?�?              �?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?      �?              �?      �?�������?333333�?      �?      �?              �?      �?                      �?      �?              �?        �>�>��?؂-؂-�?ffffff�?333333�?�������?<<<<<<�?�rO#,��?|a���?      �?      �?      �?        ZZZZZZ�?�������?              �?�������?�?              �?ffffff�?333333�?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        t�E]t�?��.���?p�}��?�Gp��?�q�q�?�q�q�?�������?�������?              �?�$I�$I�?۶m۶m�?333333�?�������?              �?      �?              �?      �?      �?                      �?              �?              �?r�q��?�q�q�?�������?UUUUUU�?              �?      �?                      �?5M�4M��?�eY�eY�?      �?        	�=����?�i��F�?F]t�E�?]t�E�?h/�����?�Kh/��?�$I�$I�?�m۶m��?              �?      �?                      �?�?<<<<<<�?      �?      �?      �?      �?              �?      �?                      �?      �?        ��8��8�?�q�q�?UUUUUU�?UUUUUU�?      �?        �����F�?W�+�ɵ?�������?UUUUUU�?ffffff�?�������?UUUUUU�?UUUUUU�?      �?              �?        ��Moz��?Y�B��?      �?              �?      �?              �?�������?�?      �?        �������?UUUUUU�?      �?      �?�������?�������?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        T:�g *�?kq�w��?��y��y�?1�0��?              �?�������?UUUUUU�?              �?      �?        �{a���?a����?������?p>�cp�?              �?�q�q�?9��8���?      �?              �?      �?�������?�������?      �?                      �?              �?�������?�������?;�;��?;�;��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        �Q�&��?�\Ų���?�������?�?�k(����?�k(���?�{a���?5�rO#,�?A��)A�?pX���o�?�?�?              �?      �?      �?      �?                      �?^Cy�5�?Q^Cy��?1�0��?��y��y�?�q�q�?r�q��?              �?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?                      �?              �?      �?        �?�?              �?UUUUUU�?�������?      �?                      �?      �?        �8��8��?9��8���?/�袋.�?F]t�E�?              �?      �?        �$I�$I�?�m۶m��?�������?�������?              �?      �?              �?      �?      �?                      �?�i��F�?GX�i���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?      �?        �袋.��?]t�E�?      �?        ;�;��?ى�؉��?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        �:��1�?�?�9�?�q�q�?r�q��?]t�E�?t�E]t�?      �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        �z�G��?{�G�z�?�.�袋�?F]t�E�?      �?        ]t�E�?F]t�E�?      �?      �?      �?                      �?�{����?�B!��?      �?      �?	�%����?h/�����?O��N���?;�;��?�?�?      �?              �?      �?      �?        �؉�؉�?;�;��?]t�E�?F]t�E�?      �?              �?              �?        ��U����?�������?333333�?ffffff�?UUUUUU�?UUUUUU�?      �?                      �?
������?��9A��?־a���?��)A��?�q�q�?�q�q�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��7��M�?d!Y�B�?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        KKKKKK�?�������?|���?|���?|��{���?���?ffffff�?333333�?      �?              �?      �?      �?                      �?�q�q�?�q�q�?      �?      �?�����?z�z��?��N��N�?�؉�؉�?]t�E]�?F]t�E�?ffffff�?333333�?      �?              �?      �?�$I�$I�?۶m۶m�?�������?333333�?      �?              �?                      �?p>�cp�?������?���k(�?(�����?      �?        �������?UUUUUU�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?              �?              �?                      �?;�;��?ى�؉��?UUUUUU�?�������?              �?      �?              �?        ZZZZZZ�?�������?      �?        �$I�$I�?۶m۶m�?�������?333333�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�
HyhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                  x#J@��ϙLq�?�           8�@              o                    �?ʲ�y��?�           �@               f                    @r�q?�?w             h@                                   @(��a��?m            �e@                                   L@�nkK�?-            @Q@                                 �A@0�,���?+            �P@       ������������������������       �                     G@               	                   �C@�����?             5@        ������������������������       �                     �?        
                           �?P���Q�?             4@                                   �?@4և���?	             ,@        ������������������������       �                      @                                  @F@�8��8��?             (@                                   �?z�G�z�?             @        ������������������������       �                      @                                  �E@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               G                    �?�E��
��?@             Z@              F                    @���@M^�?'             O@              E                    @d��0u��?&             N@              0                 �̌@�^���U�?%            �L@              /                    @���!pc�?            �@@              *                 ��@$��m��?             :@                                s@���N8�?             5@        ������������������������       �                     @                %                 ���@�q�q�?
             .@        !       "                    �?z�G�z�?             @        ������������������������       �                      @        #       $                 �|Y:@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        &       '                 ���@ףp=
�?             $@        ������������������������       �                     @        (       )                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        +       ,                    4@z�G�z�?             @        ������������������������       �                     @        -       .                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        1       2                    �?r�q��?             8@        ������������������������       �                     @        3       >                    �?�G��l��?             5@       4       5                    �?      �?	             (@        ������������������������       �                     �?        6       =                 ��&@"pc�
�?             &@       7       8                    9@ףp=
�?             $@       ������������������������       �                     @        9       :                 �?�@z�G�z�?             @        ������������������������       �                     @        ;       <                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ?       D                    ,@�����H�?             "@        @       A                    �?      �?             @        ������������������������       �                      @        B       C                 `f7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        H       _                 `f�;@և���X�?             E@       I       ^                    �?^������?            �A@       J       Y                    �?�!���?             A@       K       R                    .@�4�����?             ?@       L       Q                   �3@X�Cc�?	             ,@        M       N                 `f�)@����X�?             @        ������������������������       �                     @        O       P                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        S       X                    �?�IєX�?             1@       T       U                    �?      �?             0@       ������������������������       �                     @        V       W                 03�1@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        Z       [                   �"@�q�q�?             @        ������������������������       �                     �?        \       ]                 �|�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        `       e                    @؇���X�?             @       a       b                    @      �?             @        ������������������������       �                     �?        c       d                 ��T?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        g       h                    @�d�����?
             3@        ������������������������       �                     @        i       n                   �0@�q�q�?             (@       j       m                    @      �?              @       k       l                    @؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        p       �                 pF�,@������?           0z@       q       �                    �?$�q-�?�            q@        r       y                    8@������?             A@        s       t                 ���@�q�q�?             "@        ������������������������       �                      @        u       v                    -@և���X�?             @        ������������������������       �                      @        w       x                   �2@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        z       �                    �?HP�s��?             9@       {       |                 ���@�8��8��?             8@        ������������������������       �                     "@        }       �                 �|�=@�r����?             .@       ~                        �|=@z�G�z�?             $@        ������������������������       �                      @        �       �                   @@      �?              @       ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?X�aC�U�?�            �m@       �       �                 ��]@�;hѓ�?�            @l@        ������������������������       �        2            �S@        �       �                   �@��<D�m�?[            `b@        �       �                    >@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                   �?@`�q�0ܴ?X            �a@       �       �                   �3@���J��??            �Y@        �       �                   �2@�IєX�?             1@       ������������������������       �                     &@        �       �                 0S5 @r�q��?             @       �       �                 �?�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                   �'@`��>�ϗ?2            @U@       ������������������������       �        *            �R@        �       �                 �|�<@�C��2(�?             &@        ������������������������       �                     @        �       �                 �|�=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@��-�=��?            �C@        �       �                   @C@X�<ݚ�?             "@       �       �                    A@�q�q�?             @        ������������������������       �      �?             @        ������������������������       �                      @        �       �                   �C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     >@        �       �                   �4@�	j*D�?	             *@        �       �                    �?�q�q�?             @        �       �                  s�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    &@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    0@��[.K�?d            @b@        �       �                    �?��}*_��?             ;@       ������������������������       �        	             ,@        �       �                 X�lA@�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @        �       �                   �R@؇���X�?U            �]@       �       �                    �?(2��R�?T            �]@       �       �                    �?�z�6�?0             O@        �       �                    H@      �?             0@       �       �                 `f�A@���Q��?             $@       �       �                      @      �?              @       �       �                  �>@���Q��?             @       �       �                 X�,@@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�3Ea�$�?$             G@       �       �                   �J@"pc�
�?"             F@       �       �                 `fF:@������?             >@        ������������������������       �        
             &@        �       �                   �G@D�n�3�?             3@       �       �                 �T!@@������?             .@        �       �                   @>@�q�q�?             @       �       �                 �|Y=@      �?             @        ������������������������       �                     �?        �       �                 `fF<@�q�q�?             @       �       �                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     ,@        �       �                 03C7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @�h����?$             L@        �       �                    �?8�Z$���?             *@       �       �                   �C@z�G�z�?             $@       �       �                 ���7@�q�q�?             @        ������������������������       �                     @        �       �                   �;@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �? qP��B�?            �E@       ������������������������       �                     @@        �       �                    @�C��2(�?	             &@        �       �                  �v6@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �                           @�-���?>             Y@       �       �                    �?��[�p�?;            �W@       �       �                    �?��2(&�?             F@       ������������������������       �                     <@        �       �                    �?      �?             0@        ������������������������       �                     @        �       �                 ��UO@���Q��?             $@        ������������������������       �                      @        �       �                 0��U@      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                 �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                  �? �o_��?             I@                                 �?r�q��?             2@       ������������������������       �                     ,@                                 �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                 @     ��?             @@                                �?�z�G��?             >@       ������������������������       �        	             1@        	      
                ��#@�	j*D�?             *@        ������������������������       �                      @                              `�iJ@"pc�
�?             &@        ������������������������       �                     �?                                �B@ףp=
�?             $@        ������������������������       �                     @                                �D@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������Ӭ����?�X�>��?����<��?֖�~���?�������?�����*�?y&>�?���"��?d!Y�B�?�Mozӛ�?g��1��?Ez�rv�?              �?�a�a�?=��<���?      �?        �������?ffffff�?�$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?              �?      �?        ��؉���?;�;��?�c�1��?�s�9��?wwwwww�?DDDDDD�?:��,���?c:��,��?t�E]t�?F]t�E�?vb'vb'�?�N��N��?��y��y�?�a�a�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?�$I�$I�?۶m۶m�?              �?      �?        �������?�������?      �?              �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?        ��y��y�?1�0��?      �?      �?              �?/�袋.�?F]t�E�?�������?�������?      �?        �������?�������?      �?              �?      �?              �?      �?                      �?�q�q�?�q�q�?      �?      �?              �?      �?      �?              �?      �?                      �?              �?      �?        ۶m۶m�?�$I�$I�?_�_��?uPuP�?�������?�������?��RJ)��?���Zk��?%I�$I��?�m۶m��?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �?�?      �?      �?              �?F]t�E�?]t�E�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        Cy�5��?y�5���?      �?        �������?�������?      �?      �?۶m۶m�?�$I�$I�?              �?      �?              �?                      �?e�\x�U�?�=�S�?�؉�؉�?;�;��?xxxxxx�?�?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?                      �?q=
ףp�?{�G�z�?UUUUUU�?UUUUUU�?      �?        �������?�?�������?�������?      �?              �?      �?333333�?�������?      �?              �?              �?        ���hB�?Tn�wp٫?R��Ź�?�:Fq�c�?      �?        ��S�r
�?և���X�?      �?      �?      �?                      �?��F}g��?W�+�ɥ?______�?�?�?�?      �?        �������?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�?      �?        ]t�E�?F]t�E�?      �?        �������?�������?              �?      �?        }˷|˷�?�A�A�?r�q��?�q�q�?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        vb'vb'�?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        Q�B�
�?�z��ի�?_B{	�%�?B{	�%��?      �?        �؉�؉�?ى�؉��?              �?      �?        ۶m۶m�?�$I�$I�?=�"h8��?'u_[�?J)��RJ�?�Zk����?      �?      �?333333�?�������?      �?      �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ����7��?��,d!�?/�袋.�?F]t�E�?wwwwww�?�?      �?        l(�����?(������?wwwwww�?�?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?      �?                      �?      �?              �?      �?              �?      �?        �$I�$I�?۶m۶m�?;�;��?;�;��?�������?�������?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?              �?        ��}A�?�}A_З?      �?        ]t�E�?F]t�E�?      �?      �?      �?              �?      �?              �?      �?              �?                      �?�p=
ף�?�G�z��?m�w6�;�?�
br1�?t�E]t�?��.���?              �?      �?      �?              �?333333�?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?      �?              �?      �?              �?        �Q����?
ףp=
�?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?      �?333333�?ffffff�?              �?vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?              �?�������?�������?      �?        �������?�������?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���]hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMIhjh))��}�(h,h/h0MI��h2h3h4hph<�h=Kub������       ,                   �0@�����?�           8�@                                   �?���Q��?3             T@                               P��+@$��m��?             J@        ������������������������       �                     $@                                   @և���X�?             E@        ������������������������       �                     @                                    @^H���+�?            �B@        ������������������������       �                     2@        	                        ��T?@�����?             3@       
                        `f7@      �?             0@                                  �?���|���?             &@                                  �?      �?              @                               03�-@r�q��?             @                                 �-@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               %                    $@      �?             <@                                  �;@�ՙ/�?             5@                                  �?$�q-�?	             *@                                   @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                      @        !       "                    �?      �?              @        ������������������������       �                     @        #       $                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        &       +                    �?؇���X�?             @       '       (                    �?      �?             @        ������������������������       �                     �?        )       *                 �̌!@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        -       �                     @\��J���?�           ��@        .       �                  x#J@������?�             r@       /       ^                     �?�R�!�u�?}             i@        0       ]                    �?p�ݯ��?*             S@       1       \                    �?L�qA��?)            �R@       2       U                  �>@ޚ)�?(             R@       3       T                    �?z�):���?             I@       4       ;                    �?z�J��?            �G@        5       6                    �?�q�q�?             (@        ������������������������       �                      @        7       8                 ��";@�z�G��?             $@        ������������������������       �                     @        9       :                   �<@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        <       S                    R@�xGZ���?            �A@       =       >                 `V�9@4���C�?            �@@        ������������������������       �                     @        ?       R                    N@��
ц��?             :@       @       I                 �|�?@�z�G��?             4@        A       B                    <@և���X�?             @        ������������������������       �                     �?        C       D                 `fF<@�q�q�?             @        ������������������������       �                     @        E       H                   @>@�q�q�?             @       F       G                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        J       K                    �?8�Z$���?             *@        ������������������������       �                     @        L       Q                   �J@�<ݚ�?             "@       M       P                   `G@      �?              @       N       O                 `f�;@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        V       [                    �?�C��2(�?             6@        W       Z                 �DhF@8�Z$���?             *@       X       Y                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     �?        _       n                    �?X�'����?S             _@        `       i                    �?և���X�?
             ,@       a       h                 pf�,@�<ݚ�?             "@       b       g                    �?      �?              @       c       d                   �(@z�G�z�?             @        ������������������������       �                      @        e       f                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        j       m                    �?z�G�z�?             @        k       l                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        o       �                    �?2t3����?I            �[@       p       {                    �?U��
�??            @W@        q       z                   �J@4?,R��?             B@       r       u                   �;@(N:!���?            �A@        s       t                   �6@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        v       w                   �7@h�����?             <@       ������������������������       �                     8@        x       y                   �E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        |       �                   �A@l�b�G��?'            �L@       }       �                 `fF)@������?            �B@       ~       �                    �?�X�<ݺ?             2@              �                    5@      �?             0@        �       �                   �2@r�q��?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �        	             $@        ������������������������       �                      @        �       �                    �?�S����?             3@       �       �                   �3@d}h���?	             ,@       �       �                 �|Y;@�θ�?             *@        ������������������������       �                     @        �       �                 �|�=@�q�q�?             "@        ������������������������       �                      @        �       �                    @@؇���X�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        �       �                    �?�IєX�?
             1@        ������������������������       �                     $@        �       �                   �:@؇���X�?             @       ������������������������       �                     @        �       �                   @A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @H@f.i��n�?9            �V@       �       �                    �?������?,             Q@       �       �                 �|�=@�z�6�?(             O@        �       �                    �?�LQ�1	�?             7@       ������������������������       �        
             (@        �       �                    �?���!pc�?             &@       �       �                   �9@      �?              @        ������������������������       �                     @        �       �                 Ъb@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @T@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�ݜ�?            �C@       ������������������������       �                     >@        �       �                   @B@X�<ݚ�?             "@        ������������������������       �                     @        �       �                 8�<Q@r�q��?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 @�pX@�eP*L��?             6@       �       �                    �?���!pc�?             &@       �       �                   @J@�����H�?             "@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?"pc�
�?             &@        ������������������������       �                     �?        �       �                    �?ףp=
�?             $@       ������������������������       �                     @        �       �                 `f�h@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���@�<dVo�?�            Pu@        ������������������������       �                     ?@        �       H                  �C@xG�"��?�            `s@       �       G                   �?R�͖2�?�            �q@       �       �                    �?��e�K�?�            �p@        �       �                   @C@ҐϿ<��?)            �N@       �       �                    @8^s]e�?'             M@       �       �                    �?��N`.�?%            �K@        �       �                    �?؇���X�?             5@       �       �                    �?��S�ۿ?             .@       �       �                    �?$�q-�?	             *@        ������������������������       �                     @        �       �                 �|Y8@ףp=
�?             $@        ������������������������       �                     �?        �       �                 ���@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �@�ʻ����?             A@        �       �                   �2@"pc�
�?             &@        ������������������������       �                     �?        �       �                    �?ףp=
�?             $@       �       �                 �|�;@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �9@\X��t�?             7@       �       �                 @33"@r�q��?	             (@        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                    �?�q�q�?             @       �       �                    4@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���!pc�?             &@       �       �                    �?�q�q�?             @       �       �                    ;@      �?             @        ������������������������       �                     �?        �       �                 ��� @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       @                   �?�`�=	�?�            �i@       �       /                  �>@      �?}             h@       �                         @4@ w���?o            �d@        �       �                 �&�@�d�����?             3@        ������������������������       �                     �?        �       �                 @3�@�<ݚ�?             2@        ������������������������       �                     @        �                       0S5 @���|���?             &@       �                          �3@�q�q�?             @       �       �                   �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                �5@,N�_� �?`            �b@        ������������������������       �                     *@              .                   �?�>����?Y            �`@                                �?6uH���?P             _@                                �6@�����H�?             ;@        ������������������������       �                     �?        	                        �+@$�q-�?             :@       
                      ���@`2U0*��?             9@        ������������������������       �                     (@                              �|=@$�q-�?             *@        ������������������������       �                     @                              �|�=@�����H�?             "@                               @@      �?              @       ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                              ���@,���$�??            @X@        ������������������������       �                     �?                                 �?      �?>             X@        ������������������������       �                     .@                              ��) @�>����?2            @T@                             �|Y=@ �.�?Ƞ?#             N@       ������������������������       �                     =@                               sW@�g�y��?             ?@                              pf�@؇���X�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     8@               -                �|�=@���N8�?             5@       !      &                @3�!@z�G�z�?             4@        "      #                �|Y<@      �?             @        ������������������������       �                     �?        $      %                pf� @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        '      (                  �<@      �?             0@        ������������������������       �                     @        )      ,                   (@�����H�?             "@        *      +                ���"@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             &@        0      1                  �?@��H�}�?             9@        ������������������������       �                     @        2      3                   �?���N8�?             5@        ������������������������       �                     @        4      ?                   �?�E��ӭ�?             2@       5      <                  @@@     ��?
             0@        6      ;                d�6@@և���X�?             @       7      :                ��I @�q�q�?             @       8      9                �?�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        =      >                @3�@�<ݚ�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        A      F                8#�1@����X�?	             ,@       B      E                   �?և���X�?             @       C      D                  �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             3@        ������������������������       �                     8@        �*       h�h))��}�(h,h/h0MIKK��h2h3h4hVh<�h=Kub�����������������?��܍��?�������?333333�?vb'vb'�?�N��N��?              �?۶m۶m�?�$I�$I�?      �?        �g�`�|�?L�Ϻ��?              �?Q^Cy��?^Cy�5�?      �?      �?]t�E]�?F]t�E�?      �?      �?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�a�a�?�<��<��?;�;��?�؉�؉�?F]t�E�?]t�E�?              �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?        �.k���?���)o�?8���?�<�p�?�G�z�?ףp=
��?^Cy�5�?Cy�5��?t�@��?�K~���?9��8���?��8��8�?H�z�G�?q=
ףp�?AL� &W�?}g���Q�?�������?�������?      �?        333333�?ffffff�?              �?333333�?�������?      �?                      �?�_�_�?�A�A�?m��&�l�?'�l��&�?      �?        �؉�؉�?�;�;�?333333�?ffffff�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?;�;��?;�;��?              �?�q�q�?9��8���?      �?      �?      �?      �?              �?      �?                      �?      �?              �?                      �?      �?        ]t�E�?F]t�E�?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?        �c�1��?t�9�s�?۶m۶m�?�$I�$I�?�q�q�?9��8���?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?�������?      �?      �?              �?      �?              �?        *A��)�?�}��7��?��O?���?X`��?r�q��?�8��8��?�A�A�?|�W|�W�?۶m۶m�?�$I�$I�?              �?      �?        �$I�$I�?�m۶m��?              �?      �?      �?              �?      �?              �?        �Gp��?p�}��?��g�`��?к����?��8��8�?�q�q�?      �?      �?�������?UUUUUU�?      �?              �?      �?      �?              �?        (������?^Cy�5�?I�$I�$�?۶m۶m�?ى�؉��?�؉�؉�?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?        �?�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        �>�>��?�`�`�?�?xxxxxx�?�Zk����?J)��RJ�?d!Y�B�?Nozӛ��?              �?F]t�E�?t�E]t�?      �?      �?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �i�i�?\��[���?              �?r�q��?�q�q�?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?      �?                      �?t�E]t�?]t�E�?t�E]t�?F]t�E�?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?        /�袋.�?F]t�E�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �y�g��?�f�a��?      �?        ������?=���?̒r@d�?�ϴ5�n�?~�fߥ��?�2A�L�?mާ�d�?������?	�=����?|a���?� O	��?��oX���?�$I�$I�?۶m۶m�?�?�������?;�;��?�؉�؉�?              �?�������?�������?              �?�q�q�?�q�q�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        <<<<<<�?�������?F]t�E�?/�袋.�?      �?        �������?�������?UUUUUU�?�������?              �?      �?                      �?!Y�B�?��Moz��?�������?UUUUUU�?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?      �?        t�E]t�?F]t�E�?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?              �?      �?                      �?      �?        ��6���?�H%�e�?      �?      �?W��1 �?E���w��?Cy�5��?y�5���?              �?9��8���?�q�q�?      �?        ]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?      �?              �?        h�`�|��?���L�?      �?        �Kh/��?h/�����?k���Zk�?��RJ)��?�q�q�?�q�q�?              �?�؉�؉�?;�;��?���Q��?{�G�z�?      �?        �؉�؉�?;�;��?      �?        �q�q�?�q�q�?      �?      �?�������?�������?      �?              �?                      �?�,O"Ӱ�?���fy�?              �?      �?      �?      �?        �Kh/��?h/�����?wwwwww�?�?      �?        ��{���?�B!��?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?        �a�a�?��y��y�?�������?�������?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?      �?                      �?      �?        {�G�z�?
ףp=
�?              �?�a�a�?��y��y�?      �?        �q�q�?r�q��?      �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?9��8���?�q�q�?      �?      �?      �?              �?        �m۶m��?�$I�$I�?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?              �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�;hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       \                    �?��l�Qf�?�           8�@                                    @�������?�            �p@                                  �?BӀN��?[            �b@                                03�=@`���i��?             F@                                   D@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     D@        	                           6@88��M�?=            �Z@        
                          �2@R�}e�.�?             :@                                  �?R���Q�?             4@                                 �9@     ��?	             0@        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     @                                   ?@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        0            @T@               /                    �?\X��t�?I            �\@                                    �?���!pc�?            �K@                               �|Y8@l��\��?             A@        ������������������������       �                     @                                ���@ �Cc}�?             <@                                �Y�@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                                   �?�nkK�?             7@       ������������������������       �        
             1@                                   �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        !       .                    �?և���X�?
             5@       "       )                 �|Y=@�t����?             1@        #       $                 ���,@���Q��?             @        ������������������������       �                     �?        %       (                 `�@1@      �?             @       &       '                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        *       -                    �?r�q��?             (@        +       ,                 X��B@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        0       S                 `f7@�q�q�?,             N@       1       R                    �?��6���?             E@       2       C                   �9@      �?             C@       3       @                    �?�ՙ/�?             5@       4       ?                   �7@�q�q�?             2@       5       <                    �?���Q��?
             .@       6       ;                 pff@�q�q�?             (@       7       :                    4@����X�?             @        8       9                 P��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        =       >                 �!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        A       B                     @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        D       Q                    �?ҳ�wY;�?             1@       E       L                    �?     ��?             0@       F       G                 �|�;@X�<ݚ�?             "@        ������������������������       �                     @        H       I                 �|�=@�q�q�?             @        ������������������������       �                     @        J       K                    A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        M       P                   �0@؇���X�?             @       N       O                 �|�;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       W                    �?�����H�?             2@        U       V                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        X       Y                 ��T?@@4և���?
             ,@        ������������������������       �                      @        Z       [                    %@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ]       h                    *@R�����?           �{@        ^       _                     @�X����?             6@        ������������������������       �                      @        `       a                    �?      �?	             ,@        ������������������������       �                     @        b       e                    �?���|���?             &@        c       d                 ��!>@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        f       g                 03�8@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        i       �                 `ff:@�����?           pz@       j       u                     @�\���?�            ps@        k       l                 `f�)@ ������?)            �O@        ������������������������       �                     >@        m       t                    �?Pa�	�?            �@@       n       o                   @D@���7�?             6@       ������������������������       �                     .@        p       s                    ,@؇���X�?             @        q       r                   �F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        v       �                    �?��a�n`�?�             o@       w       �                    �?�TG!u�?�            �n@        x       �                  �v6@$G$n��?+            �R@       y       �                    �?0�й���?*            @R@       z       �                    �?�LQ�1	�?)            @Q@       {       �                 �|Y=@�r����?"             N@        |       �                    �?���Q��?             $@       }       �                 ��=@      �?              @       ~                        ��y@z�G�z�?             @        ������������������������       �                     �?        �       �                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|�=@`2U0*��?             I@       �       �                    �?P���Q�?             D@        ������������������������       �                     .@        �       �                 ���@HP�s��?             9@        ������������������������       �                     @        �       �                 ��(@�����H�?
             2@       ������������������������       ��r����?             .@        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?�����H�?             "@       ������������������������       �                     @        �       �                 ��y&@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��|�N
�?u            �e@       �       �                   �7@������?c             b@        �       �                 @3�@`2U0*��?!             I@       ������������������������       �                     9@        �       �                 pf� @HP�s��?             9@        �       �                   �1@�q�q�?             @        ������������������������       �                      @        �       �                   �4@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �        
             3@        �       �                    �?�W�{�5�?B            �W@       �       �                 �?�@$�3c�s�?A            �W@       �       �                   �8@ �q�q�?!             H@        �       �                 `fF@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �F@        �       �                   �;@�3Ea�$�?              G@        �       �                 pf� @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 @3�@r�q��?             E@        �       �                   �?@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �A@      �?              @       ������������������������       ����Q��?             @        ������������������������       ��q�q�?             @        �       �                 ��) @�FVQ&�?            �@@        ������������������������       �                     0@        �       �                 ��y @�t����?             1@        ������������������������       �                     �?        �       �                 �|�=@      �?             0@       ������������������������       �                     &@        �       �                    ?@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 pf� @h�����?             <@        �       �                 P�@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     �?        �       �                   �<@      �?E             \@        �       �                     �?�5��?             ;@       �       �                    �?j���� �?             1@       �       �                   �8@�eP*L��?             &@        ������������������������       �                     @        �       �                   �;@؇���X�?             @       ������������������������       �                     @        �       �                 `f�D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        �       �                 �nc@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                  "&d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �9@ףp=
�?             $@       ������������������������       �                     @        �       �                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?z�G�z�?3            @U@       �       �                    �?�w��@�?'            �O@       �       �                      @�q�q��?             H@       �       �                  �?@� ��1�?            �D@        �       �                    @@D�n�3�?             3@        �       �                 �|�=@�<ݚ�?             "@       �       �                    <@      �?              @        ������������������������       �                     @        �       �                 ��2>@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �F@���Q��?             $@        ������������������������       �                     @        �       �                   @Q@�q�q�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                   �=@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        �       �                 �|�>@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                     �?�q�q�?             .@       �       �                   �E@�n_Y�K�?	             *@       �       �                  x#J@�q�q�?             @        ������������������������       �                     �?        �       �                   �B@z�G�z�?             @        �       �                 `f�K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �H@؇���X�?             @        �       �                   �G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �                          �?���7�?             6@                               pU�t@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������}<����?�/���?��9����?\�qA��?ـl@6 �?�7���M�?F]t�E�?F]t�E�?      �?      �?              �?      �?                      �?����f��?+J�#��?�;�;�?'vb'vb�?333333�?333333�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?��Moz��?!Y�B�?t�E]t�?F]t�E�?�������?------�?              �?۶m۶m�?%I�$I��?�������?333333�?              �?      �?        d!Y�B�?�Mozӛ�?              �?UUUUUU�?�������?      �?                      �?�$I�$I�?۶m۶m�?�������?�������?�������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?UUUUUU�?�m۶m��?�$I�$I�?              �?      �?              �?                      �?�������?�������?=��<���?b�a��?      �?      �?�<��<��?�a�a�?UUUUUU�?UUUUUU�?333333�?�������?�������?�������?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?�q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?�������?      �?                      �?              �?      �?                      �?�q�q�?�q�q�?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?      �?        �������?UUUUUU�?              �?      �?        �'�R0�?9a��>��?]t�E]�?�E]t��?              �?      �?      �?              �?]t�E]�?F]t�E�?�������?333333�?              �?      �?        �������?UUUUUU�?              �?      �?        4F���?��/�	�?�F�zm�?
���*��?��}��}�?AA�?      �?        |���?|���?�.�袋�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �s�9��?�c�1Ƹ?@�O%��?�����߸?к����?���L�?����?����Ǐ�?��Moz��?Y�B��?�������?�?�������?333333�?      �?      �?�������?�������?      �?              �?      �?              �?      �?                      �?              �?���Q��?{�G�z�?ffffff�?�������?      �?        q=
ףp�?{�G�z�?      �?        �q�q�?�q�q�?�������?�?      �?              �?        �q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?fGi�?+���}��?��y�!�?C:o1��?���Q��?{�G�z�?      �?        q=
ףp�?{�G�z�?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        �ĩ�sK�?Fڱa��?1���\A�?x6�;��?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        ����7��?��,d!�?      �?      �?      �?                      �?�������?UUUUUU�?�q�q�?r�q��?              �?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?>����?|���?      �?        <<<<<<�?�?              �?      �?      �?      �?        �������?�������?              �?      �?              �?        �m۶m��?�$I�$I�?]t�E�?F]t�E�?      �?                      �?      �?              �?              �?      �?h/�����?/�����?ZZZZZZ�?�������?]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�}��}��?AA�?�������?UUUUUU�?������?������?l(�����?(������?9��8���?�q�q�?      �?      �?      �?        333333�?�������?              �?      �?              �?        �������?333333�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?      �?                      �?              �?      �?        �$I�$I�?۶m۶m�?      �?                      �?UUUUUU�?UUUUUU�?;�;��?ى�؉��?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �.�袋�?F]t�E�?۶m۶m�?�$I�$I�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ� �thG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       H                     �?���*1�?�           8�@                                   �?gO�~k�?l            @d@                                   �?j�g�y�?+             O@                                  �?#z�i��?            �D@        ������������������������       �                     2@                                �;|r@�û��|�?             7@                                  �?�q�q�?             5@                                  H@     ��?             0@       	       
                    9@�eP*L��?             &@        ������������������������       �                      @                                �|�;@X�<ݚ�?             "@        ������������������������       �                      @                                   C@և���X�?             @                               �|�=@�q�q�?             @                               ��2>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                  �B@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                   �?���N8�?             5@                                 �4@$�q-�?
             *@                                   �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @                =                    �?���o_�?A             Y@       !       "                    �?:W��S��?1             S@        ������������������������       �                     �?        #       $                    �?�EH,���?0            �R@        ������������������������       �                     4@        %       <                    �?�2�o�U�?#            �K@       &       1                  i?@l��
I��?"             K@        '       (                 ��$:@�ՙ/�?             5@        ������������������������       �                     @        )       0                 `fF<@�r����?	             .@       *       +                 03k:@"pc�
�?             &@        ������������������������       �                      @        ,       -                 �|�?@�<ݚ�?             "@        ������������������������       �                     �?        .       /                   �J@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        2       3                  x#J@�C��2(�?            �@@       ������������������������       �                     3@        4       ;                 03�M@d}h���?             ,@        5       6                    9@      �?             @        ������������������������       �                     �?        7       :                 `f�K@���Q��?             @       8       9                   �C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        >       G                    �?r�q��?             8@       ?       B                    �?z�G�z�?             4@       @       A                    �?�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @        C       F                 ���R@؇���X�?             @        D       E                   @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        I       h                     @L [ܝ�?W           (�@        J       a                    �?nN[]�?`            �c@       K       L                    �?Ҿ ؞��?D            �[@        ������������������������       �                     @        M       R                    �?�B�����?@             Z@        N       O                   �B@��S�ۿ?             >@       ������������������������       �                     3@        P       Q                    D@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        S       `                    �?xL��N�?,            �R@       T       U                    �?����˵�?$            �M@        ������������������������       �                      @        V       Y                    4@�}�+r��?#            �L@        W       X                    &@�<ݚ�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        Z       [                   @D@@��8��?             H@       ������������������������       �                     ?@        \       _                   �*@�IєX�?	             1@       ]       ^                   @G@�����H�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     .@        b       c                   �8@z�G�z�?            �F@        ������������������������       �                     (@        d       e                    �?���!pc�?            �@@       ������������������������       �                     4@        f       g                    ,@�	j*D�?
             *@        ������������������������       �                     @        ������������������������       �                     "@        i       �                    �?�]��NH�?�            �x@        j       �                   �B@���3L�?E             [@       k       �                    �? U����?>            �X@        l       w                    4@�*/�8V�?            �G@        m       r                    �?��S���?             .@        n       o                    �?z�G�z�?             @        ������������������������       �                     @        p       q                 ��!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        s       t                 �*@���Q��?             $@        ������������������������       �                      @        u       v                    @      �?              @        ������������������������       �                      @        ������������������������       �                     @        x       �                 �|�=@     ��?             @@       y       ~                 �|Y<@r�q��?             >@        z       }                    �?      �?	             0@       {       |                 P�@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     @               �                    '@d}h���?
             ,@       �       �                 ���@8�Z$���?	             *@        �       �                 �Y�@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���4@��B����?!             J@       �       �                 ��.@^������?            �A@        �       �                    �?     ��?
             0@       �       �                   �1@X�Cc�?	             ,@        �       �                    �?r�q��?             @       �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�S����?             3@        ������������������������       �                     @        �       �                 �|�7@d}h���?             ,@        ������������������������       �                     �?        �       �                    @@8�Z$���?             *@       �       �                 ��1@      �?              @        ������������������������       �                     @        �       �                 03C3@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @������?             1@        �       �                    @���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�8��8��?	             (@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     "@        �       �                    #@�r����?�            �q@        �       �                 @3�4@�q�q�?             8@       ������������������������       �                     ,@        ������������������������       �                     $@        �       �                   �<@���(`�?�            Pp@        �       �                    �?�}�+r��?D            �\@        �       �                    �?���!pc�?             &@       �       �                    5@����X�?             @        ������������������������       �                     @        �       �                   �6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��&@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �9@ f^8���?>            �Y@       �       �                 �?�@�d���?3            �U@        ������������������������       �                     F@        �       �                   �4@ �#�Ѵ�?            �E@       �       �                    �?@4և���?             <@       �       �                    �?�����?             5@       �       �                   �2@�}�+r��?             3@        �       �                 pf� @r�q��?             @        �       �                    1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        �       �                    2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        �       �                 0�@@      �?             0@       ������������������������       �        	             ,@        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y=@�q��/��?a            `b@        �       �                    �?      �?             $@       �       �                    �?      �?              @        ������������������������       �                     @        �       �                 ���"@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?���	���?Z             a@        �       �                    �?�t����?             1@       �       �                 �|�=@      �?             0@       �       �                 ���@ףp=
�?	             $@        ������������������������       �                     @        �       �                    �?r�q��?             @       �       �                   @@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�.�?�P�?K             ^@        �       �                    �?���}<S�?             7@       �       �                 X��A@�����?             5@       �       �                   `3@�KM�]�?             3@       ������������������������       �                     0@        �       �                 03�7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �                          �?�$��y��?<            @X@       �                         �C@ą%�E�?7            @V@       �                       ��C@��UV�?,            �Q@       �       �                 pf�@t�e�í�?+            �P@        ������������������������       �        	             1@        �                          �?ףp=
�?"             I@       �                          @C@�����H�?            �F@       �       �                   @@@@4և���?             E@       �       �                   �@     ��?             @@        �       �                 �|Y>@�q�q�?             @        ������������������������       �                     �?        �       �                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�=@XB���?             =@       �       �                 ��) @�nkK�?             7@       ������������������������       �                     3@        �       �                 �̜!@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������`l����??'��d�?��"e���?�n���?��{���?B!�B�?ە�]���?�+Q��?              �?8��Moz�?��,d!�?UUUUUU�?UUUUUU�?      �?      �?t�E]t�?]t�E�?      �?        �q�q�?r�q��?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?        333333�?�������?              �?      �?                      �?�a�a�?��y��y�?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?              �?��Q���?=
ףp=�?����k�?���k(�?      �?        7�i�6�?�_,�Œ�?              �?־a��?�S�<%��?Lh/����?h/�����?�a�a�?�<��<��?      �?        �?�������?F]t�E�?/�袋.�?              �?�q�q�?9��8���?      �?              �?      �?              �?      �?                      �?]t�E�?F]t�E�?      �?        I�$I�$�?۶m۶m�?      �?      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?UUUUUU�?�������?�������?�������?�؉�؉�?ى�؉��?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �? n�D�?��#��w�?�A�A�?˷|˷|�?q��$�?��2���?      �?        b'vb'v�?;�;��?�?�������?              �?F]t�E�?/�袋.�?      �?                      �?>�S��?L�Ϻ��?W'u_�?��/���?      �?        �5��P�?(�����?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?        �?�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?              �?              �?        �������?�������?              �?t�E]t�?F]t�E�?              �?vb'vb'�?;�;��?              �?      �?        ��q����?���H�?&���^B�?�%���^�?A�_)P��?`)P�W
�?AL� &W�?�٨�l��?�������?�?�������?�������?              �?      �?      �?      �?                      �?333333�?�������?              �?      �?      �?              �?      �?              �?      �?UUUUUU�?�������?      �?      �?UUUUUU�?�������?              �?      �?                      �?۶m۶m�?I�$I�$�?;�;��?;�;��?      �?      �?              �?      �?                      �?      �?                      �?O��N���?ى�؉��?_�_��?uPuP�?      �?      �?%I�$I��?�m۶m��?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?^Cy�5�?(������?              �?۶m۶m�?I�$I�$�?      �?        ;�;��?;�;��?      �?      �?              �?      �?      �?      �?                      �?              �?xxxxxx�?�?�������?333333�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?        �������?�?�������?�������?              �?      �?        g��o��?Ȥx�L��?�5��P�?(�����?F]t�E�?t�E]t�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?H%�e�?��VCӝ?�:���C�?Ȥx�L��?      �?        �/����?�}A_Ч?n۶m۶�?�$I�$I�?=��<���?�a�a�?�5��P�?(�����?�������?UUUUUU�?      �?      �?      �?                      �?      �?              �?              �?      �?      �?                      �?      �?              �?              �?      �?      �?              �?      �?              �?      �?        /����?և���X�?      �?      �?      �?      �?              �?333333�?�������?      �?                      �?      �?        V��,���?P�9��J�?<<<<<<�?�?      �?      �?�������?�������?      �?        �������?UUUUUU�?�������?�������?      �?      �?      �?              �?              �?                      �?�?wwwwww�?ӛ���7�?d!Y�B�?=��<���?�a�a�?�k(���?(�����?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ����?W?���?�as���?��g<�?2~�ԓ��?6��9�?�1����?�rv��?      �?        �������?�������?�q�q�?�q�q�?n۶m۶�?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?GX�i���?�{a���?�Mozӛ�?d!Y�B�?      �?              �?      �?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��1hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       j                     @�,�٧��?�           8�@                                   )@0Z� ���?�            ps@                                  �F@r�q��?             B@                                  �?ףp=
�?             >@        ������������������������       �                     �?                                   �? 	��p�?             =@        ������������������������       �                      @        ������������������������       �                     ;@        	       
                   �J@      �?             @        ������������������������       �                     @        ������������������������       �                     @               %                    �?���Q��?�            0q@                                   @�Z]]Y�?S            �`@                                ��1V@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               $                 03�<@���7�?Q            �`@               #                    �?ףp=
�?"             N@              "                 ���;@�r����?            �F@                                   �?@4և���?             E@        ������������������������       �                     @                                  �2@�8��8��?             B@                                  :@P���Q�?             4@        ������������������������       �                     �?        ������������������������       �        
             3@               !                   �E@      �?	             0@                                  �?��S�ۿ?             .@        ������������������������       �                      @                                   �7@$�q-�?             *@                                   �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             .@        ������������������������       �        /             R@        &       ?                    �?6�|�3�?[            �a@        '       8                    �?R���Q�?             D@       (       7                   �H@�q�q�?             8@       )       6                     �?p�ݯ��?             3@       *       +                   �7@     ��?             0@        ������������������������       �                      @        ,       5                    C@X�Cc�?	             ,@       -       4                 �̾w@      �?             (@       .       3                 �|Y<@"pc�
�?             &@       /       0                   �9@�q�q�?             @        ������������������������       �                     @        1       2                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        9       >                     �?      �?             0@       :       =                    �?�<ݚ�?             "@       ;       <                 p"�X@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        @       A                    $@��%3�?B            @Y@        ������������������������       �                     $@        B       M                 ��$:@��0%�?<            �V@        C       L                   @A@l��\��?             A@        D       E                 �|�<@@�0�!��?             1@       ������������������������       �                     $@        F       K                   �3@և���X�?             @       G       H                 �|�=@      �?             @        ������������������������       �                      @        I       J                    @@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     1@        N       i                 03�M@��h!��?"            �L@       O       h                     �?�q�q�?             H@       P       _                    �?���|���?             F@       Q       ^                    K@�q�q�?             >@       R       ]                 ��yC@�G��l��?             5@       S       T                 �|�<@      �?             0@        ������������������������       �                     @        U       \                   �H@�eP*L��?	             &@       V       W                 03k:@      �?              @        ������������������������       �                     �?        X       [                   �>@؇���X�?             @        Y       Z                 `f�<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        `       a                  x#J@և���X�?             ,@        ������������������������       �                     @        b       c                    7@�q�q�?             "@        ������������������������       �                     �?        d       e                    A@      �?              @        ������������������������       �                     @        f       g                   �C@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        k       �                    �?&S��:�?�             y@        l       }                 03@6C�z��?E            �\@        m       |                    �?t�F�}�?             �I@       n       o                    �? �o_��?             I@        ������������������������       �                     "@        p       q                   �6@,���i�?            �D@        ������������������������       �                      @        r       {                    �?$�q-�?            �C@       s       t                   �<@�L���?            �B@        ������������������������       �                     @        u       v                    �?ףp=
�?             >@        ������������������������       �                     (@        w       x                  s�@r�q��?             2@        ������������������������       �                     @        y       z                 �|Y=@�θ�?	             *@        ������������������������       �                     �?        ������������������������       �r�q��?             (@        ������������������������       �                      @        ������������������������       �                     �?        ~       �                 03�:@�q�q�?%            �O@              �                    �?      �?              L@       �       �                    �?(N:!���?            �A@       �       �                 P��+@���y4F�?	             3@        ������������������������       �                     @        �       �                   �-@����X�?             ,@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 X��B@"pc�
�?             &@       �       �                    �?ףp=
�?             $@        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     0@        �       �                    �?�G��l��?             5@       �       �                    �?      �?
             (@       �       �                 �&�)@ףp=
�?	             $@        �       �                 �|�4@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @"pc�
�?�            �q@        �       �                 ���A@��<b���?             7@       �       �                    @ףp=
�?             4@        �       �                    �?�q�q�?             @        ������������������������       �                      @        �       �                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                     @        �       �                    �?���B��?�            pp@       �       �                    �?���9yw�?�            �m@        �       �                 ��}@��c:�?             G@        ������������������������       �                     @        �       �                    �?X�Cc�?             E@       �       �                    �?\�Uo��?             C@       �       �                    �?�q�q�?             8@       �       �                  �#@8����?             7@       �       �                   �@r�q��?
             2@        �       �                   �A@      �?              @       �       �                    4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                 �[$@z�G�z�?             @        ������������������������       �                     @        �       �                 ��&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�<@      �?	             ,@       �       �                    4@����X�?             @        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���.@����X�?             @        ������������������������       �                     �?        �       �                 �|Y>@r�q��?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �?�@X��R9�?x             h@        �       �                    �?��V�I��?:            �W@       �       �                   �7@X;��?7            @V@        ������������������������       �                     ?@        �       �                   �8@�8���?$             M@        �       �                 `fF@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��@ 7���B�?!             K@        ������������������������       �                     7@        �       �                 �|�=@`Jj��?             ?@       �       �                 �|Y=@      �?             0@        ������������������������       �                     @        �       �                  sW@"pc�
�?	             &@        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                     @        �       �                 @3�@�����H�?>            �X@        �       �                   �9@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �?@      �?              @        ������������������������       �                     �?        �       �                   �A@և���X�?             @       ������������������������       ��q�q�?             @        ������������������������       �      �?             @        �       �                    �?����\�?7            �V@       �       �                    �? wVX(6�?1            @T@       �       �                 �|�=@�n���?*             R@       �       �                   �2@���U�?             �L@        �       �                 ��Y @r�q��?             (@        �       �                    1@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                    �F@        �       �                   �?@z�G�z�?
             .@        �       �                 �̌!@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        �       �                    5@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        �       �                    @ �q�q�?             8@       �       �                 ��l&@�X�<ݺ?             2@        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������&��jq�?:�g *�?AW o��?_��oH��?�������?UUUUUU�?�������?�������?              �?������?�{a���?              �?      �?              �?      �?              �?      �?        �������?333333�?z�rv��?�՘HT�?      �?      �?              �?      �?        F]t�E�?�.�袋�?�������?�������?�?�������?�$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?�������?ffffff�?      �?                      �?      �?      �?�?�������?              �?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?      �?              �?                      �?              �?�k:`�?E�)͋?�?�������?�������?�������?�������?^Cy�5�?Cy�5��?      �?      �?              �?%I�$I��?�m۶m��?      �?      �?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?      �?              �?              �?      �?9��8���?�q�q�?      �?      �?              �?      �?              �?              �?        :5r���?���Q`�?              �?�Q�Q�?�������?------�?�������?ZZZZZZ�?�������?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?              �?      �?      �?              �?        Hp�}�?p�}��?UUUUUU�?UUUUUU�?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?1�0��?��y��y�?      �?      �?              �?t�E]t�?]t�E�?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?              �?        �$I�$I�?۶m۶m�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?      �?      �?                      �?      �?              �?        \���(\�?H�z�G�?~��G�?��Gp�?777777�?�������?
ףp=
�?�Q����?              �?�����?8��18�?              �?�؉�؉�?;�;��?}���g�?L�Ϻ��?      �?        �������?�������?      �?        �������?UUUUUU�?      �?        ى�؉��?�؉�؉�?              �?�������?UUUUUU�?      �?              �?        UUUUUU�?UUUUUU�?      �?      �?�A�A�?|�W|�W�?(������?6��P^C�?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?/�袋.�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?��y��y�?1�0��?      �?      �?�������?�������?�������?�������?              �?      �?              �?                      �?�q�q�?�q�q�?              �?      �?              �?        /�袋.�?F]t�E�?��Moz��?��,d!�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?        �X�J���?��2�*��?��Y��?���s��?-d!Y��?�7��Mo�?              �?%I�$I��?�m۶m��?�5��P^�?6��P^C�?UUUUUU�?UUUUUU�?d!Y�B�?8��Moz�?�������?UUUUUU�?      �?      �?      �?      �?      �?                      �?      �?              �?        �������?�������?              �?      �?      �?      �?                      �?              �?      �?      �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        BN�­�?��葲?<�����?AL� &W�?�u�{���?�E(B�?      �?        j��FX�?a���{�?      �?      �?              �?      �?        	�%����?h/�����?      �?        ���{��?�B!��?      �?      �?      �?        /�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?              �?              �?        �q�q�?�q�q�?r�q��?�q�q�?      �?              �?      �?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?.؂-؂�?�>�>�?k~X�<�?�<ݚ�?r�q��?r�qǱ?	�#����?p�}��?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        �������?�������?      �?      �?      �?                      �?      �?        9��8���?�q�q�?      �?              �?      �?              �?      �?              �?        �������?UUUUUU�?��8��8�?�q�q�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�JIhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       
                   @���*1�?�           8�@              S                    �?~ @���?�           ��@                                    @���f)w�?�            �l@                                  �?H�Swe�?S            @_@                                   �?�>����?4            @T@       ������������������������       �        !             J@                                   B@V�a�� �?             =@              	                 ��Y)@      �?             8@        ������������������������       �                     &@        
                           �?�θ�?
             *@        ������������������������       �                     @                                   <@      �?              @                                  �7@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                   �?���Q��?             @                                 �'@      �?             @                                 �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     F@               N                   @B@��WV��?@             Z@              K                    @,�[I'��?9            �W@              ,                    �?F�����?6            �V@               '                    �?r�q��?             >@                               �|Y8@�����H�?             2@        ������������������������       �                     @               "                  ��@8�Z$���?
             *@                !                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        #       $                 ���@�C��2(�?             &@        ������������������������       �                     �?        %       &                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        (       +                 ��.@      �?
             (@        )       *                   �-@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        -       F                 03�1@�������?             N@       .       A                    �?j���� �?            �I@       /       <                  �#@X�<ݚ�?             B@       0       9                   �7@X�<ݚ�?             ;@       1       8                    �?X�<ݚ�?	             2@       2       3                 ���@��.k���?             1@        ������������������������       �                      @        4       5                    4@�����H�?             "@        ������������������������       �                     @        6       7                 pff@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        :       ;                 �|Y>@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        =       @                 ��&@�����H�?             "@       >       ?                    4@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        B       C                    4@�q�q�?             .@        ������������������������       �                     @        D       E                   �.@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        G       H                    �?�����H�?             "@        ������������������������       �                     @        I       J                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        L       M                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        O       R                   @C@ףp=
�?             $@        P       Q                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        T       W                    ,@��늓��?           �|@        U       V                    @�IєX�?             1@       ������������������������       �        
             0@        ������������������������       �                     �?        X       �                     �?��>܀�?           �{@        Y       x                    �?��:��?7            @V@        Z       q                    �?j���� �?             A@       [       j                 ��UO@�z�G��?             4@       \       i                    �?z�G�z�?
             .@       ]       ^                 `f&;@���!pc�?             &@        ������������������������       �                     �?        _       `                 ���<@z�G�z�?             $@        ������������������������       �                     @        a       h                 p�i@@����X�?             @       b       g                   �H@      �?             @       c       d                 ��2>@�q�q�?             @        ������������������������       �                     �?        e       f                  �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        k       p                    �?���Q��?             @       l       m                 0c@      �?             @        ������������������������       �                      @        n       o                 X�l@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        r       w                   �H@և���X�?             ,@       s       t                 �UcV@���!pc�?             &@       ������������������������       �                     @        u       v                 Ј�V@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        y       �                  i?@\�����?"            �K@        z       �                    K@      �?             8@       {       |                 �̌*@�X����?             6@        ������������������������       �                     @        }       �                 �|Y=@���y4F�?	             3@        ~                          @>@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 `fF<@@4և���?             ,@       �       �                   @G@z�G�z�?             @        �       �                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        �       �                    �?f���M�?             ?@       �       �                   �A@� �	��?             9@        ������������������������       �                     @        �       �                    H@�G��l��?             5@       �       �                    �?X�<ݚ�?             2@        �       �                 ��yC@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    7@�eP*L��?             &@        ������������������������       �                      @        �       �                 03�M@X�<ݚ�?             "@       �       �                    A@����X�?             @        ������������������������       �                     @        �       �                  x#J@      �?             @        ������������������������       �                     �?        �       �                 `�iJ@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�(̶h�?�            @v@       �       �                 0��D@h�ƄbB�?�            Pr@       �       �                   �3@�����H�?�             r@        �       �                     @�d�����?             C@        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        �       �                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �2@��R[s�?            �A@       �       �                   �1@�X����?             6@       �       �                   �0@������?             .@       �       �                 pFD!@�q�q�?             (@       �       �                 pf�@      �?              @        ������������������������       �                     @        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��@և���X�?             @        ������������������������       �                      @        �       �                 ��Y @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 0S5 @8�Z$���?             *@       �       �                 �?�@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 @3�@h�N?���?�            @o@       �       �                    ?@      �?O             `@       �       �                 �|Y=@�$��y��?@            @X@       �       �                    �?8�Z$���?!             J@        �       �                   �<@�eP*L��?             &@       �       �                 ��y@����X�?             @        ������������������������       �                      @        �       �                 ���@���Q��?             @        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���@������?            �D@        �       �                 ���@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �A@        �       �                 �|�=@����?�?            �F@       �       �                 �Y�@ qP��B�?            �E@        �       �                    �?ףp=
�?	             $@       �       �                 ���@      �?              @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                    �@@        ������������������������       �                      @        �       �                   @@@��a�n`�?             ?@        ������������������������       �                     @        �       �                 �?�@�����H�?             ;@       ������������������������       �                     8@        ������������������������       �                     @        �       �                 ��q1@�.ߴ#�?H            �^@       �       �                     @��?^�k�?@            @Z@        �       �                 �|�=@ qP��B�?            �E@        �       �                   �'@�����H�?             "@        ������������������������       �                      @        �       �                    �?؇���X�?             @        ������������������������       �                      @        �       �                 �|Y<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     A@        �       �                 �|�=@�g�y��?)             O@       ������������������������       �                    �D@        �       �                 ��)"@�����?             5@       ������������������������       �                     0@        �       �                    (@���Q��?             @       �       �                   �?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �4@@�0�!��?             1@        ������������������������       �                     @        ������������������������       �                     ,@        �       �                    ;@���Q��?             @        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       	                   �?$Q�q�?)            �O@       �       �                    �?�NW���?!            �J@        �       �                 03�-@      �?              @        ������������������������       �                     @        �       �                 �|�=@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �                            @`Ӹ����?            �F@        ������������������������       �                     ,@                                 �?`Jj��?             ?@        ������������������������       �                     @                                 5@HP�s��?             9@                                 �?�<ݚ�?             "@                                �2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        ������������������������       �                     $@        ������������������������       �                     4@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������`l����??'��d�?HO.�7s�?pa���?��G���?��λ�?�~j�t��?X9��v�?h/�����?�Kh/��?              �?a���{�?��{a�?      �?      �?              �?�؉�؉�?ى�؉��?              �?      �?      �?      �?      �?      �?                      �?              �?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?��N��N�?��؉���?�
br1�?���F}g�?؂-؂-�?�>�>��?UUUUUU�?�������?�q�q�?�q�q�?              �?;�;��?;�;��?      �?      �?              �?      �?        F]t�E�?]t�E�?              �?�������?�������?              �?      �?              �?      �?      �?      �?      �?                      �?              �?�������?�������?ZZZZZZ�?�������?�q�q�?r�q��?r�q��?�q�q�?�q�q�?r�q��?�?�������?              �?�q�q�?�q�q�?      �?        �������?UUUUUU�?              �?      �?                      �?9��8���?�q�q�?      �?                      �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?r�q��?�q�q�?      �?                      �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �������?�������?      �?      �?      �?                      �?      �?        ��e�:}�?T,h�?�?�?              �?      �?        ���Od�?g�$��o�?�x�3��?�as���?�������?ZZZZZZ�?ffffff�?333333�?�������?�������?F]t�E�?t�E]t�?              �?�������?�������?      �?        �m۶m��?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?              �?        �������?333333�?      �?      �?              �?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?t�E]t�?F]t�E�?              �?      �?      �?      �?                      �?      �?        ߰�k��?A��)A�?      �?      �?]t�E]�?�E]t��?      �?        (������?6��P^C�?333333�?�������?      �?                      �?�$I�$I�?n۶m۶�?�������?�������?      �?      �?              �?      �?                      �?              �?      �?        ��RJ)��?��Zk���?�Q����?)\���(�?      �?        ��y��y�?1�0��?r�q��?�q�q�?�$I�$I�?۶m۶m�?              �?      �?        t�E]t�?]t�E�?      �?        �q�q�?r�q��?�$I�$I�?�m۶m��?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �JV����?��MmjS�?4!RzdI�?d�n-ܴ�?�q�q�?�q�q�?Cy�5��?y�5���?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        X|�W|��?PuPu�?�E]t��?]t�E]�?wwwwww�?�?UUUUUU�?UUUUUU�?      �?      �?      �?        �������?�������?      �?              �?        �$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?        ;�;��?;�;��?�m۶m��?�$I�$I�?      �?                      �?      �?        �v��/�?�I+��?      �?      �?����?W?���?;�;��?;�;��?]t�E�?t�E]t�?�m۶m��?�$I�$I�?      �?        333333�?�������?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?p>�cp�?������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��I��I�?l�l��?��}A�?�}A_З?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?        �c�1��?�s�9��?              �?�q�q�?�q�q�?      �?                      �?�K�`m�?XG��).�?_�_��?�A�A�?��}A�?�}A_З?�q�q�?�q�q�?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?      �?        ��{���?�B!��?      �?        =��<���?�a�a�?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ZZZZZZ�?�������?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ~��}���?AA�?萚`���?�x+�R�?      �?      �?      �?        333333�?�������?              �?      �?        ?�>��?l�l��?      �?        ���{��?�B!��?      �?        q=
ףp�?{�G�z�?9��8���?�q�q�?      �?      �?      �?                      �?      �?              �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��NhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       L                     �?���%&�?�           8�@               +                  x#J@o����?o            �e@               *                    �?�#��ؒ�?-            @Q@              )                    �?     ��?+             P@                                  �?¦	^_�?*             O@                                  �H@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        	                           �?�T`�[k�?%            �J@        
                        �ܵ<@�θ�?	             *@        ������������������������       �                      @                                `f�A@���!pc�?             &@                                  �?�q�q�?             "@                                �>@և���X�?             @                                Y>@�q�q�?             @                               X��E@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                `fF:@R���Q�?             D@        ������������������������       �                     "@               (                   @J@¦	^_�?             ?@              '                   �H@և���X�?             5@              &                   �F@p�ݯ��?             3@              %                 `f�D@      �?
             ,@              $                   @>@���|���?             &@              #                 `fF<@      �?              @              "                 �|�?@�q�q�?             @                !                 �|�<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     @        ,       -                    �?� ���?B            @Z@       ������������������������       �        )            �P@        .       =                    �?      �?             C@       /       6                 p"�X@
;&����?             7@       0       5                    I@�	j*D�?	             *@       1       4                   �8@ףp=
�?             $@        2       3                 ���Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        7       <                    �?�z�G��?             $@       8       ;                   @E@      �?             @       9       :                   �:@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        >       K                    @��S���?             .@       ?       @                 `�iJ@      �?
             ,@        ������������������������       �                      @        A       J                 03�U@�q�q�?	             (@       B       I                 `��T@�z�G��?             $@       C       D                    �?      �?              @        ������������������������       �                     �?        E       H                    <@����X�?             @        F       G                    7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        M       b                    /@6�����?X           Ȁ@        N       [                    @8^s]e�?)             M@       O       Z                 ��3@@4և���?             E@        P       W                    �?r�q��?             2@       Q       R                 P��+@r�q��?             (@       ������������������������       �                     @        S       V                    �?���Q��?             @       T       U                   �-@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        X       Y                 ���2@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     8@        \       ]                    �?      �?             0@        ������������������������       �                     @        ^       a                    @�����H�?             "@        _       `                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        c       �                    �?@O'D��?/           �}@       d       �                    �?��
�d8�?�            py@        e       n                    �?U��
�?9            @W@        f       g                 ���@ܷ��?��?             =@        ������������������������       �                      @        h       i                    �? 7���B�?             ;@       ������������������������       �        
             3@        j       m                    �?      �?              @        k       l                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        o       x                  ��@     ��?'             P@        p       w                    �?�FVQ&�?            �@@       q       r                 ���@ףp=
�?             4@       ������������������������       �                     (@        s       t                 �|=@      �?              @        ������������������������       �                      @        u       v                 �|�=@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     *@        y       �                    �?��a�n`�?             ?@       z       �                    �?�+$�jP�?             ;@       {       |                 �|Y=@��<b���?             7@        ������������������������       �                     @        }       ~                     @ףp=
�?             4@        ������������������������       �                      @               �                 �|Y?@�����H�?             2@       �       �                    �?8�Z$���?	             *@        ������������������������       �                      @        ������������������������       �"pc�
�?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                  �v6@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?��ۭ���?�            �s@       �       �                     @�}���?�            0s@        �       �                    �?6�}0S��?@            �[@        �       �                    �?z�G�z�?             >@       �       �                 `f&'@�X�<ݺ?             2@        �       �                   �J@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             *@        �       �                   �7@�q�q�?             (@        ������������������������       �                      @        �       �                   �E@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?*             T@       �       �                   @A@�[|x��?#            �O@       �       �                 �|Y=@X�EQ]N�?            �E@       �       �                    &@(;L]n�?             >@        �       �                    5@ףp=
�?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �        	             4@        �       �                   �'@�	j*D�?	             *@       ������������������������       �                     @        �       �                 �|�=@�q�q�?             @        ������������������������       �                     @        �       �                    @@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     4@        ������������������������       �                     1@        �       �                 ��) @���G�?�            �h@       �       �                    �?���	���?Y             a@       �       �                    ;@�[|x��?S            �_@        �       �                   �9@�y��*�?#             M@       �       �                 �?$@ �h�7W�?             �J@        �       �                   �2@ȵHPS!�?             :@        �       �                 P��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �5@���}<S�?             7@        ������������������������       �                     "@        �       �                    �?؇���X�?             ,@        �       �                    8@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     ;@        �       �                 @3�@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �&B@ =[y��?0             Q@        ������������������������       �                     8@        �       �                 �Yu@t��ճC�?              F@        ������������������������       �                     �?        �       �                    �? �#�Ѵ�?            �E@        ������������������������       �                     �?        �       �                   �>@���N8�?             E@       ������������������������       �                     9@        �       �                 @3�@�t����?             1@       �       �                   �?@z�G�z�?             $@        ������������������������       �                     �?        �       �                 �?�@�����H�?             "@        ������������������������       �                     @        �       �                   �A@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                   �4@���!pc�?             &@        �       �                 03�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    9@�������?'             N@        �       �                 Ь�#@�nkK�?             7@       ������������������������       �                     3@        �       �                    �?      �?             @        �       �                 �[$@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��!@^H���+�?            �B@        �       �                    �?�n_Y�K�?             *@        ������������������������       �                     @        �       �                 �|�>@      �?             $@        �       �                 pf� @����X�?             @        ������������������������       �                     @        �       �                 �|Y<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���.@�q�q�?             8@        ������������������������       �                      @        �       �                    �?     ��?             0@       �       �                 �T�C@�z�G��?             $@        ������������������������       �                      @        �       �                 �|�>@      �?              @       �       �                    ;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                 ��1@      �?             @       �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     @b�2�tk�?1             R@        �       �                    �?�X����?             6@       ������������������������       �        
             .@        ������������������������       �                     @        �                          �?�-���?              I@        �       �                    5@      �?             (@        ������������������������       �                      @        �                          �?ףp=
�?             $@       �       �                 �|Y=@؇���X�?             @        ������������������������       �                     @        �                         S�2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?�KM�]�?             C@                             03c"@r�q��?             8@                              �|Y7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?              	                   �?�����?             5@        ������������������������       �                     @        
                          @�����H�?             2@                             ��T?@"pc�
�?             &@                               �>@ףp=
�?             $@       ������������������������       �                     @                                �A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             ,@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������g *��?�0���M�?5�rO#,�?�FX�i�?F��Q�g�?s��\;0�?      �?      �?��Zk���?�RJ)���?UUUUUU�?UUUUUU�?              �?      �?        ���!5��?"5�x+��?ى�؉��?�؉�؉�?      �?        F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?              �?        �������?�������?      �?        ��Zk���?�RJ)���?�$I�$I�?۶m۶m�?^Cy�5�?Cy�5��?      �?      �?F]t�E�?]t�E]�?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?              �?                      �?      �?                      �?              �?�r)�r)�?Z�5Z�5�?              �?      �?      �?�Mozӛ�?Y�B��?;�;��?vb'vb'�?�������?�������?      �?      �?              �?      �?                      �?      �?        ffffff�?333333�?      �?      �?      �?      �?      �?                      �?      �?              �?        �?�������?      �?      �?              �?�������?�������?ffffff�?333333�?      �?      �?              �?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?              �?                      �?      �?        �*��o��?1��� ��?	�=����?|a���?�$I�$I�?n۶m۶�?UUUUUU�?�������?UUUUUU�?�������?              �?�������?333333�?      �?      �?      �?                      �?              �?UUUUUU�?�������?              �?      �?                      �?      �?      �?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        v=���?(
�o���?@v\�_��?�&�����?��O?���?X`��?a���{�?��=���?      �?        h/�����?	�%����?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?     ��?      �?>����?|���?�������?�������?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?              �?        �c�1��?�s�9��?/�����?B{	�%��?��,d!�?��Moz��?              �?�������?�������?      �?        �q�q�?�q�q�?;�;��?;�;��?      �?        /�袋.�?F]t�E�?      �?              �?              �?      �?      �?                      �?�?m�K�?�Kz���?aD���)�?}9Y�?��yJ��?߰�k��?�������?�������?�q�q�?��8��8�?�������?�������?              �?      �?                      �?�������?�������?      �?        333333�?ffffff�?              �?      �?              �?      �?]�u]�u�?EQEQ�?w�qG�?qG�wĽ?�������?�?�������?�������?      �?      �?      �?              �?        vb'vb'�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?        �~=��?����?V��,���?P�9��J�?]�u]�u�?EQEQ�?�4�rO#�?GX�i��?��sHM0�?"5�x+��?��N��N�?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?        ӛ���7�?d!Y�B�?      �?        ۶m۶m�?�$I�$I�?333333�?�������?              �?      �?              �?              �?        �������?�������?              �?      �?        �������?�������?      �?        �E]t��?t�E]t�?              �?�/����?�}A_Ч?      �?        ��y��y�?�a�a�?      �?        <<<<<<�?�?�������?�������?              �?�q�q�?�q�q�?      �?        �������?�������?      �?              �?      �?      �?        F]t�E�?t�E]t�?      �?      �?      �?                      �?      �?        �������?�������?�Mozӛ�?d!Y�B�?      �?              �?      �?      �?      �?              �?      �?              �?        L�Ϻ��?�g�`�|�?ى�؉��?;�;��?              �?      �?      �?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?              �?        UUUUUU�?�������?      �?              �?      �?ffffff�?333333�?      �?              �?      �?�������?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        �8��8��?9��8���?]t�E]�?�E]t��?              �?      �?        �G�z��?�p=
ף�?      �?      �?      �?        �������?�������?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�k(���?(�����?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        =��<���?�a�a�?      �?        �q�q�?�q�q�?/�袋.�?F]t�E�?�������?�������?      �?              �?      �?              �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ2�3hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K煔h2h3h4hph<�h=Kub��������       �                 03[L@�����?�           8�@              S                    �?B�=�o��?~           �@               6                    �?�T
Z��?p            �d@                                   @*��)^�?W             `@                                  �E@     ��?)             P@                                 �;@`'�J�?"            �I@                                   �?�����?             5@        ������������������������       �                     "@        	       
                   �9@r�q��?             (@       ������������������������       �                     "@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     >@                                   �?�	j*D�?             *@                                  �?z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @                                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               %                 �|�<@�n_Y�K�?.            @P@                                  @�ʻ����?             A@        ������������������������       �                     @               $                    �?��X��?             <@              !                    �?��H�}�?             9@                                 �5@և���X�?
             ,@        ������������������������       �                     @                                   �7@�q�q�?             "@                               pff@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        "       #                 P�@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        &       5                   @D@�n`���?             ?@       '       4                 03�7@r�q��?             >@       (       )                    �? �Cc}�?             <@       ������������������������       �        
             0@        *       -                    �?      �?             (@        +       ,                 �|�=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        .       3                     @�����H�?             "@       /       0                 03�1@      �?              @       ������������������������       �                     @        1       2                 03C3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        7       R                    @��+��?            �B@       8       O                 ��p@@)O���?             B@       9       :                 ��Y@�q�q�?             ;@        ������������������������       �                      @        ;       H                    �? �o_��?             9@       <       E                 �|Y=@r�q��?
             (@       =       >                     @ףp=
�?             $@        ������������������������       �                     @        ?       D                    @r�q��?             @       @       C                    1@z�G�z�?             @        A       B                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        F       G                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       N                   @C@�n_Y�K�?             *@       J       M                    *@z�G�z�?             $@        K       L                 ��T?@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        P       Q                     @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        T       [                    @�)���?           �{@        U       X                    �?����X�?             5@        V       W                    @�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        Y       Z                    �?�q�q�?             (@        ������������������������       �                     @        ������������������������       �                     @        \       �                   �R@�Ǣ3F�?           `z@       ]       �                 ��D:@�<����?           0z@       ^       u                    �?H����?�            Pu@        _       r                    �?d}h���?             E@       `       o                    �?:�&���?            �C@       a       l                 83�0@<���D�?            �@@       b       c                 ���@@4և���?             <@        ������������������������       �        	             ,@        d       e                   �5@؇���X�?
             ,@        ������������������������       �                     �?        f       g                     @$�q-�?	             *@        ������������������������       �                     @        h       i                 �|�:@ףp=
�?             $@        ������������������������       �                      @        j       k                   @@      �?              @        ������������������������       �      �?             @        ������������������������       �                     @        m       n                   �2@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        p       q                 �&�)@      �?             @        ������������������������       �                     @        ������������������������       �                     @        s       t                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        v       �                    �?`5�#�t�?�            �r@       w       x                    )@h�Y���?�            Pr@        ������������������������       �                     �?        y       z                    �?F��}��?�            @r@        ������������������������       �                     ;@        {       |                 �?�@V^���?�            �p@        ������������������������       �        =            @X@        }       �                    �?�����?^             e@       ~       �                   �<@$��$�L�?W            �c@               �                    �?�IєX�?$             Q@       �       �                     @�i�y�?!            �O@        ������������������������       �                     :@        �       �                 0S5 @@-�_ .�?            �B@        �       �                    3@����X�?             @        �       �                    1@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     >@        �       �                     @���Q��?             @        ������������������������       �                     �?        �       �                 pf(@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    $@�r����?3            �V@        �       �                   �"@���"͏�?            �B@       �       �                 @3�@��a�n`�?             ?@        �       �                   �A@      �?             (@       ������������������������       �      �?              @        ������������������������       �      �?             @        ������������������������       �                     3@        ������������������������       �                     @        �       �                     @ �h�7W�?            �J@       �       �                 �|�=@t��ճC�?             F@        �       �                    1@؇���X�?             @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �@@@-�_ .�?            �B@        ������������������������       �                     *@        �       �                   @A@�8��8��?             8@        �       �                    1@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        �       �                   @D@P���Q�?             4@        ������������������������       �                     $@        �       �                    �?ףp=
�?             $@       �       �                   �F@�����H�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     $@        ������������������������       �                     @        �       �                  �>@��Sݭg�?4            �S@        �       �                    �?)O���?             B@       �       �                    �?�f7�z�?             =@       �       �                    K@$��m��?             :@       �       �                   `G@�KM�]�?             3@       �       �                   �F@"pc�
�?	             &@       �       �                 ��";@ףp=
�?             $@        ������������������������       �                     @        �       �                 �ܵ<@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                  x#J@@4և���?             E@       ������������������������       �                     @@        �       �                 `�iJ@�z�G��?             $@        ������������������������       �                     �?        �       �                 �|�>@�<ݚ�?             "@       �       �                   �;@؇���X�?             @        �       �                    7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                      @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @@�0�!��?=            �Y@       �       �                    �?�*v��?9            @X@       �       �                    "@��?^�k�?(            �Q@        ������������������������       �                      @        ������������������������       �        '             Q@        �       �                    �?�5��?             ;@       �       �                 ���Q@�t����?
             1@        ������������������������       �                     @        �       �                    �?�eP*L��?             &@       �       �                   �G@      �?              @       �       �                 p�w@����X�?             @       �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 03�U@���Q��?             $@       �       �                    :@r�q��?             @        ������������������������       �                     @        �       �                 03�M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                  �6f@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub������������������?��܍��?$�ՄD}�?��T�v�?��ί=��?��(��?�'�	{��?��=aO�?      �?      �?�?�������?�a�a�?=��<���?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?;�;��?vb'vb'�?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ى�؉��?;�;��?�������?<<<<<<�?              �?n۶m۶�?%I�$I��?{�G�z�?
ףp=
�?۶m۶m�?�$I�$I�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        ]t�E�?F]t�E�?              �?      �?              �?        �c�1��?�9�s��?UUUUUU�?�������?۶m۶m�?%I�$I��?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?        *�Y7�"�?�S�n�?��8��8�?9��8���?UUUUUU�?UUUUUU�?      �?        �Q����?
ףp=
�?UUUUUU�?�������?�������?�������?              �?UUUUUU�?�������?�������?�������?      �?      �?              �?      �?                      �?              �?      �?      �?      �?                      �?ى�؉��?;�;��?�������?�������?      �?      �?      �?                      �?              �?      �?        �q�q�?�q�q�?              �?      �?              �?        m��q�`�?MΡ8�}�?�$I�$I�?�m۶m��?�q�q�?�q�q�?              �?      �?        �������?�������?      �?                      �?��R��H�?&�k]���?w���|�?L����?�=��c��?�N8ᄳ?I�$I�$�?۶m۶m�?�A�A�?�o��o��?|���?|���?n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?      �?        �������?�������?      �?              �?      �?      �?      �?      �?        333333�?�������?      �?                      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?2R��;.�?���A�?�)=�$�?d�n-ܴ�?              �?��Ǐ?�?����?      �?         �{�c�?�E���?      �?        =��<���?�a�a�?��]-n��?�3���?�?�?�������?AA�?      �?        S�n0E�?к����?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?              �?        333333�?�������?      �?              �?      �?              �?      �?        �������?�?v�)�Y7�?*�Y7�"�?�s�9��?�c�1Ƹ?      �?      �?      �?      �?      �?      �?      �?                      �?��sHM0�?"5�x+��?�E]t��?t�E]t�?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        S�n0E�?к����?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?        ffffff�?�������?      �?        �������?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?              �?              �?              �?              �?        �|˷|��?�i�i�?9��8���?��8��8�?a���{�?O#,�4��?vb'vb'�?�N��N��?(�����?�k(���?F]t�E�?/�袋.�?�������?�������?              �?�������?�������?      �?                      �?      �?                      �?      �?              �?              �?        n۶m۶�?�$I�$I�?      �?        ffffff�?333333�?              �?9��8���?�q�q�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?              �?�������?ZZZZZZ�?�i�n�'�?��Id��?�A�A�?_�_��?      �?                      �?/�����?h/�����?�������?�������?              �?]t�E�?t�E]t�?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJk�ahG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������       N                    �?	dm#��?�           8�@                                   �?|��?���?�            �g@                                    @��t���?6            �S@                                0Cd=@�����?             E@                                ��@5@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �A@        	                        X�,A@����>�?            �B@       
                           �?4�2%ޑ�?            �A@                                H�%@      �?             $@        ������������������������       �                     @                                   �?����X�?             @        ������������������������       �                     @                                   �?�q�q�?             @                                  5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                   �?H%u��?             9@                               �|�9@�8��8��?             8@        ������������������������       �                     @                                ���@�����?             5@        ������������������������       �                      @        ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                      @               /                   �:@x��}�?J            �[@               ,                   �9@r�q��?             8@              !                     �?X�<ݚ�?             2@                                 ��)e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        "       +                   �6@X�Cc�?             ,@       #       *                    @      �?	             $@       $       '                    �?����X�?             @       %       &                 ��y@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        (       )                 ��}@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        -       .                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        0       9                 ��K.@"Z�l�?7            �U@       1       8                    �?@�E�x�?            �H@       2       3                     @ 7���B�?             ;@        ������������������������       �                     @        4       7                    �?�nkK�?             7@       5       6                 �|Y=@P���Q�?             4@        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     @        ������������������������       �                     6@        :       ;                 ��.@4�B��?            �B@        ������������������������       �                      @        <       M                 @��v@����X�?            �A@       =       L                    I@r٣����?            �@@       >       ?                 ��Y9@�q�q�?             8@        ������������������������       �                     @        @       K                    �?���Q��?             4@       A       J                    �?և���X�?	             ,@       B       I                     �?�n_Y�K�?             *@       C       H                   @@@�q�q�?             (@       D       E                 ���<@z�G�z�?             @        ������������������������       �                     @        F       G                 ��2>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        O       |                    �?����S��?J           P�@        P       Y                    (@����X�?g            @c@        Q       X                    �?      �?             8@       R       W                    "@؇���X�?	             ,@       S       V                    @$�q-�?             *@        T       U                 ��zT@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     $@        Z       k                     @؇>���?W            @`@       [       j                    �?����!p�?:             V@       \       i                 `fF:@�C��2(�?$            �K@       ]       h                    L@��hJ,�?             A@       ^       c                   �9@<���D�?            �@@        _       b                   �3@�q�q�?             @       `       a                   �4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        d       e                   �E@�>����?             ;@       ������������������������       �                     4@        f       g                    5@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                    �@@        l       {                 ��Y1@X�Cc�?             E@       m       z                   �:@���Q��?             9@       n       s                   �!@j���� �?             1@       o       p                   �6@X�<ݚ�?             "@        ������������������������       �                     @        q       r                   �9@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        t       y                    �?      �?              @        u       v                    4@�q�q�?             @        ������������������������       �                     �?        w       x                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             1@        }       �                 `��S@@���j�?�             w@       ~       �                     �?�D�d@6�?�            Pv@               �                   �<@      �?             H@        �       �                    �?և���X�?             @       �       �                 `f�D@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �E@� ��1�?            �D@       �       �                 �|Y>@ �o_��?             9@       �       �                    �?��S�ۿ?	             .@       �       �                   �>@@4և���?             ,@       �       �                 �|Y=@؇���X�?             @        ������������������������       �                     �?        �       �                 `fF<@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��I*@���Q��?             $@        ������������������������       �                      @        �       �                   @@@      �?              @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �H@      �?             0@        �       �                    �?      �?              @       �       �                 `f�;@r�q��?             @        �       �                 ��:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�b�E�V�?�            Ps@       �       �                 `�X#@��}����?�            �p@       �       �                     @8v�YeK�?q            �g@        ������������������������       �                     @        �       �                    7@`Jj��?m            @g@        �       �                   �2@`����֜?#            �Q@        �       �                 ��@P���Q�?	             4@        ������������������������       �                     $@        �       �                 ��Y @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     I@        �       �                   �C@�q3�M��?J             ]@       �       �                    �?d۬����??            @W@       �       �                   @C@�=C|F�?;            �U@       �       �                   @8@�̨�`<�?:            @U@        �       �                 `fF@      �?              @        �       �                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��) @�C��2(�?5            @S@       �       �                   �@�����?-            �P@        �       �                 �|�<@�8��8��?             8@        ������������������������       �                     "@        �       �                   @@@�r����?             .@       �       �                 �&B@�<ݚ�?             "@       �       �                 pf�@      �?              @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ?@ qP��B�?            �E@       ������������������������       �                     A@        �       �                   �@@�����H�?             "@       �       �                 �?�@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                 0S%"@���Q��?             $@        �       �                 X��@@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �|�=@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     7@        �       �                    �?�(�Tw�?3            �S@       �       �                    ?@ _�@�Y�?%             M@       ������������������������       �                     B@        �       �                 0��D@���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        ������������������������       �                     4@        �       �                     @���� �?            �D@        �       �                    :@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?������?             A@        ������������������������       �                     @        �       �                 `f2@�חF�P�?             ?@        �       �                    %@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @HP�s��?             9@       �       �                 ���A@ףp=
�?             4@       �       �                    �?؇���X�?	             ,@       ������������������������       �                     "@        �       �                 ��T?@���Q��?             @       �       �                    @      �?             @       �       �                    +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?���|���?             &@        �       �                    5@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������"iD��?&�-w���?{	�%���?	�%����?^-n����?�td�@T�?�a�a�?=��<���?�$I�$I�?۶m۶m�?              �?      �?                      �?���L�?�u�)�Y�?�A�A�?�������?      �?      �?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?���Q��?)\���(�?UUUUUU�?UUUUUU�?              �?�a�a�?=��<���?      �?                      �?      �?              �?        pX���o�?A��)A�?UUUUUU�?UUUUUU�?r�q��?�q�q�?      �?      �?              �?      �?        %I�$I��?�m۶m��?      �?      �?�$I�$I�?�m۶m��?�������?�������?      �?                      �?      �?      �?      �?                      �?      �?              �?        UUUUUU�?�������?              �?      �?        ʚ���)�?֔5eMY�?և���X�?9/���?	�%����?h/�����?      �?        �Mozӛ�?d!Y�B�?ffffff�?�������?              �?      �?              �?              �?        �Y7�"��?L�Ϻ��?              �?�m۶m��?�$I�$I�?>���>�?|���?UUUUUU�?UUUUUU�?      �?        333333�?�������?۶m۶m�?�$I�$I�?ى�؉��?;�;��?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?                      �?      �?              �?              �?              �?                      �?X�i���?O#,�4��?�$I�$I�?�m۶m��?      �?      �?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?      �?              �?         �����?�����?]t�E�?/�袋.�?F]t�E�?]t�E�?�������?KKKKKK�?|���?|���?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?h/�����?�Kh/��?              �?�$I�$I�?�m۶m��?              �?      �?              �?                      �?              �?%I�$I��?�m۶m��?�������?333333�?�������?ZZZZZZ�?�q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?      �?        d!Y�B�?���7��?}��|���?���й?      �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        ������?������?
ףp=
�?�Q����?�������?�?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?      �?                      �?      �?              �?        �������?333333�?      �?              �?      �?      �?      �?      �?                      �?              �?      �?      �?      �?      �?�������?UUUUUU�?      �?      �?      �?                      �?      �?              �?              �?        �jch���?��,�?��Dz�r�?��[�ը?��sK���?�a�+�?      �?        ���{��?�B!��?�������?�A�A�?ffffff�?�������?      �?        �������?�������?              �?      �?              �?        �rO#,��?�i��F�?7�p�7�?Hy�G�?�C��:��?J��/�?�������?�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ]t�E�?F]t�E�?g��1��?���@��?UUUUUU�?UUUUUU�?      �?        �������?�?9��8���?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��}A�?�}A_З?      �?        �q�q�?�q�q�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?        333333�?�������?�������?333333�?              �?      �?        �������?�������?      �?                      �?              �?      �?              �?        p��o���?�A�A�?#,�4�r�?�{a���?      �?        �.�袋�?F]t�E�?      �?                      �?      �?        jW�v%j�?,Q��+�?�$I�$I�?۶m۶m�?              �?      �?        xxxxxx�?�?              �?�Zk����?��RJ)��?      �?      �?              �?      �?        q=
ףp�?{�G�z�?�������?�������?۶m۶m�?�$I�$I�?      �?        333333�?�������?      �?      �?      �?      �?              �?      �?              �?                      �?      �?              �?        F]t�E�?]t�E]�?�������?�������?              �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ6ޤhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                    �?]@f�
�?�           8�@                                 �0@�|R���?            �}@                                   :@��Q���?             D@                                  �?�5��?             ;@                                  !@�q�q�?             8@        ������������������������       �                     @                                   �?X�<ݚ�?
             2@        ������������������������       �                     "@        	       
                 pFD!@�����H�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@               W                     @F��Á�?           0{@               $                 ��/@�5�X�k�?p            `e@               #                   @I@�1��u�?1            @R@              "                    �?���h%��?,            �O@                                  �?�̚��?*            �N@                                   :@�����H�?             2@                                  �6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  �B@��S�ۿ?             .@       ������������������������       �                     $@                                  �D@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �? �#�Ѵ�?            �E@        ������������������������       �                      @                                  �@@������?            �D@       ������������������������       �                     <@                !                   @A@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     $@        %       R                    �?Tt�ó��??            �X@       &       Q                   �M@N֩	%��?:            @V@       '       (                    7@:�1�(��?7            @U@        ������������������������       �                     @        )       2                    �?L����?4            @T@        *       1                     �?(;L]n�?             >@       +       ,                   �H@���N8�?             5@       ������������������������       �        
             .@        -       0                 ,w�U@r�q��?             @        .       /                    K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        3       N                    �?t�F�}�?"            �I@       4       M                     �?���!pc�?             F@       5       F                 `f�B@�	j*D�?            �C@       6       ?                 ���=@      �?             2@       7       :                 `f&;@�q�q�?             "@        8       9                   @D@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ;       <                 ��=@r�q��?             @        ������������������������       �                     @        =       >                 X��E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        @       A                  �>@�q�q�?             "@        ������������������������       �                     @        B       E                 X�lA@      �?             @       C       D                   �@@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        G       H                 �UP@؇���X�?             5@       ������������������������       �                     ,@        I       J                  �}S@և���X�?             @        ������������������������       �                      @        K       L                 X�,@@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        O       P                 �̾w@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        S       V                    �?�<ݚ�?             "@        T       U                   �B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        X       q                    �?�F.< �?�            �p@        Y       d                 ���@��H�}�?-            �R@        Z       c                    �?��2(&�?             6@       [       \                   �6@؇���X�?             5@        ������������������������       �                      @        ]       b                 �|�=@�}�+r��?             3@       ^       _                 �|=@�C��2(�?             &@        ������������������������       �                     @        `       a                 ���@      �?              @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        e       j                    �?��k��?            �J@        f       g                    �?��2(&�?             6@        ������������������������       �                      @        h       i                    �?R���Q�?             4@       ������������������������       �        	             1@        ������������������������       �                     @        k       p                 ��$1@�חF�P�?             ?@       l       o                    �?@4և���?             <@        m       n                 �|Y=@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             2@        ������������������������       �                     @        r       �                    �?�+$�jP�?n            �g@        s       �                 ��&@��+7��?             7@       t       �                   �"@�����?             3@       u       �                    9@z�G�z�?             .@       v                           �?      �?              @       w       x                    4@      �?             @        ������������������������       �                     �?        y       z                   �6@���Q��?             @        ������������������������       �                      @        {       ~                   �7@�q�q�?             @       |       }                 @3�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                  �#@      �?             @        ������������������������       �                      @        �       �                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�=@��Lɿ��?`            �d@       �       �                 �?$@���U�?E            �\@        �       �                 ��@H%u��?             9@       ������������������������       �                     5@        ������������������������       �      �?             @        �       �                 ��) @ }�Я��?6            @V@       ������������������������       �        $             Q@        �       �                 pf� @���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        �       �                 �&B@R�}e�.�?             J@        ������������������������       �        	             4@        �       �                   @@@     ��?             @@        �       �                 @3�@����X�?             ,@        ������������������������       �                     @        �       �                    ?@      �?              @        �       �                 �̌!@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 d�6@@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �C@�<ݚ�?             2@       �       �                 @3�@���|���?             &@        �       �                   @C@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                  x#J@�=Ϯϸ�?�            �m@       �       �                    @B&�/��?s             f@       �       �                    �?~�����?`            `b@       �       �                 ��.@�|�
��?3            @U@        �       �                     @X�<ݚ�?             "@        ������������������������       �                     �?        �       �                    �?      �?              @       �       �                    �?      �?             @       �       �                 ���,@�q�q�?             @       �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��)@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   @C@$�Z����?+             S@       �       �                    �?pH����?#            �P@       �       �                 039@�>����?             K@        �       �                    �?\-��p�?             =@       �       �                    �?@�0�!��?	             1@        ������������������������       �                      @        �       �                 ���1@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                 03�7@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     9@        �       �                   �6@�θ�?             *@       �       �                  �:@      �?             @        ������������������������       �                      @        �       �                     @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 03;@X�<ݚ�?             "@        �       �                   �E@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @G@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?t�7��?-             O@        �       �                    -@���|���?	             &@        ������������������������       �                      @        �       �                     @�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    :@L紂P�?$            �I@       �       �                    �?z�G�z�?             D@       �       �                    �?(N:!���?            �A@       �       �                    �?���7�?             6@       �       �                    5@�X�<ݺ?             2@        �       �                 �Y�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     @        �       �                     @�θ�?	             *@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    $@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                    +@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        �       �                 pfv2@r�q��?             >@        ������������������������       �                     @        �       �                    @�>����?             ;@        ������������������������       �                     &@        �       �                    @      �?             0@        ������������������������       �                     @        �       �                    @�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �                          �?0B��D�?'            �M@       �                          �?      �?             H@       �       �                   @E@l��\��?             A@       ������������������������       �                     ;@        �                       p"W@և���X�?             @                                 �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                 �?d}h���?             ,@                             �ES@����X�?             @                                @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        	                         �?z�G�z�?             @       
                         �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                  �?؇���X�?             @                              �(\�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?"pc�
�?             &@        ������������������������       �                     �?                                  �?ףp=
�?             $@                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������ߺ?9���?C����v�?&N��[��?�c�H;�?�������?333333�?/�����?h/�����?UUUUUU�?UUUUUU�?              �?�q�q�?r�q��?              �?�q�q�?�q�q�?      �?      �?      �?              �?                      �?+�_����?�%@�Z�?o"���&�?"���&��?�s�Ν;�?�1bĈ�?v]�u]��?EQEQ�??�%C���?�u�y���?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?        �?�������?              �?�������?�������?      �?                      �?�/����?�}A_Ч?      �?        p>�cp�?������?      �?        ;�;��?;�;��?              �?      �?                      �?      �?        /�����?h�����?��x�3�?s����?�������?�������?              �?�5?,R�?#e�����?�?�������?�a�a�?��y��y�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?777777�?�������?F]t�E�?t�E]t�?vb'vb'�?;�;��?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?      �?                      �?      �?        �m۶m��?�$I�$I�?      �?                      �?      �?        �q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?|��|�?>����?{�G�z�?
ףp=
�?��.���?t�E]t�?۶m۶m�?�$I�$I�?              �?�5��P�?(�����?]t�E�?F]t�E�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?        oe�Cj��?"5�x+��?t�E]t�?��.���?              �?333333�?333333�?              �?      �?        �Zk����?��RJ)��?n۶m۶�?�$I�$I�?�������?�������?              �?      �?              �?                      �?/�����?B{	�%��?Y�B��?zӛ����?^Cy�5�?Q^Cy��?�������?�������?      �?      �?      �?      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?              �?      �?      �?      �?              �?      �?              �?      �?                      �?�������?rY1P»?	�#����?p�}��?)\���(�?���Q��?      �?              �?      �?�я~���?p�\��?      �?        ��y��y�?�a�a�?              �?      �?        'vb'vb�?�;�;�?      �?              �?      �?�$I�$I�?�m۶m��?              �?      �?      �?      �?      �?      �?                      �?      �?      �?      �?                      �?9��8���?�q�q�?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        Jݗ�V�?[4��}�?�z���?�
���?K���+�?[��5;j�?�?�������?r�q��?�q�q�?              �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?              �?      �?              �?      �?        l(�����?�5��P^�?z�rv��?�1���?h/�����?�Kh/��?�{a���?a����?�������?ZZZZZZ�?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�؉�؉�?ى�؉��?      �?      �?              �?      �?      �?              �?      �?                      �?�q�q�?r�q��?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?SJ)��R�?��Zk���?]t�E]�?F]t�E�?              �?9��8���?�q�q�?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?ffffff�?ffffff�?|�W|�W�?�A�A�?�.�袋�?F]t�E�?��8��8�?�q�q�?      �?      �?      �?                      �?      �?              �?        ى�؉��?�؉�؉�?      �?      �?              �?      �?        /�袋.�?F]t�E�?              �?      �?        �������?333333�?              �?      �?              �?        �������?UUUUUU�?              �?�Kh/��?h/�����?      �?              �?      �?      �?        9��8���?�q�q�?              �?      �?        ��}ylE�?�A�I��?      �?      �?�������?------�?              �?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?        ۶m۶m�?I�$I�$�?�$I�$I�?�m۶m��?      �?      �?              �?      �?        �������?�������?      �?      �?              �?      �?                      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?/�袋.�?F]t�E�?              �?�������?�������?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��{hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       Z                    �?ʡ�;S��?�           8�@               Y                 ���Q@0,Tg��?�            �o@              T                    @�g��@(�?            @i@                                   @��nk�?t             g@                                   �?(�s���?6             U@                                  L@4և����?#             L@                                  �? �h�7W�?!            �J@                                   �?      �?              @       	       
                 03�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 ��9@`Ӹ����?            �F@       ������������������������       �                     9@                                  �E@ףp=
�?             4@       ������������������������       �        	             .@                                  @H@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     <@               S                   �>@� �	��?>             Y@              "                 ��@�û��|�?8             W@                                 s@��2(&�?             6@        ������������������������       �                     @               !                    �?@�0�!��?
             1@                               �|Y:@      �?	             0@        ������������������������       �                     @                                  ��@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        #       0                    �?��(@��?*            �Q@        $       /                 ��.@���N8�?             5@       %       .                    �?�q�q�?	             (@       &       -                    �?      �?              @       '       (                 P��+@���Q��?             @        ������������������������       �                      @        )       *                   �7@�q�q�?             @        ������������������������       �                     �?        +       ,                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        1       P                    �?և���X�?            �H@       2       3                    '@���Q��?            �F@        ������������������������       �                     @        4       G                   �*@#z�i��?            �D@       5       F                 �|�=@П[;U��?             =@       6       C                    �?�q�q�?             8@       7       B                    �?�z�G��?             4@       8       9                    3@�<ݚ�?	             2@        ������������������������       �                     �?        :       A                 @3�@@�0�!��?             1@        ;       >                 pff@�q�q�?             "@        <       =                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ?       @                   �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        D       E                   �3@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        H       O                    �?�8��8��?             (@       I       J                   �.@�����H�?             "@        ������������������������       �                     @        K       N                 03�0@r�q��?             @        L       M                 �|�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        Q       R                 @34@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        U       V                    @�X�<ݺ?             2@        ������������������������       �                     @        W       X                 ���3@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     I@        [       �                 pF�,@"~��F��?           �|@       \       ]                    ,@��X�-�?�            `q@        ������������������������       �                     �?        ^       u                 �?�@�C�gr~�?�            Pq@       _       l                    �?��
���?[            �b@        `       a                 03S@؇���X�?             5@        ������������������������       �                     �?        b       i                   @@R���Q�?             4@       c       d                   �6@�r����?	             .@        ������������������������       �                     �?        e       f                 ���@@4և���?             ,@        ������������������������       �                     @        g       h                 �|=@      �?              @        ������������������������       �                     @        ������������������������       �      �?              @        j       k                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        m       n                 ��]@�7�	|��?M             `@       ������������������������       �        3            �V@        o       t                    �?P�Lt�<�?             C@       p       s                 �Yu@�?�|�?            �B@        q       r                    :@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     A@        ������������������������       �                     �?        v       �                    �?�N̸��?H            �_@       w       z                 @3�@\#r��?D            �^@        x       y                    :@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        {       �                   `!@���^���?@            �\@        |       }                    �? �Cc}�?              L@        ������������������������       �                     �?        ~       �                 �|�=@lGts��?            �K@              �                   �:@�r����?            �F@       �       �                   �3@$�q-�?             :@       �       �                   �1@8�Z$���?             *@        ������������������������       �                     @        �       �                   �2@      �?              @        �       �                 ��Y @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 0S5 @z�G�z�?             @       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     *@        �       �                 �|Y<@���y4F�?             3@        ������������������������       �                      @        �       �                 ��) @�t����?
             1@       ������������������������       �                     ,@        �       �                 pf� @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                     @���#�İ?             �M@       �       �                   �)@ �#�Ѵ�?            �E@        ������������������������       �                     4@        �       �                    @@���}<S�?             7@        ������������������������       �                     &@        �       �                   �*@r�q��?             (@       �       �                   �A@����X�?             @        ������������������������       �                     �?        �       �                   �C@r�q��?             @        ������������������������       �                     @        �       �                    G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             0@        �       �                   �5@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     �?�"W9���?p            �f@        �       �                    @@H�z�G�?3             T@        �       �                    K@:ɨ��?            �@@       �       �                   @G@d}h���?             <@       �       �                    �?�q�q�?             2@        �       �                    �?�q�q�?             @       �       �                 �|�;@z�G�z�?             @        ������������������������       �                     �?        �       �                 X�,@@      �?             @       �       �                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @>@�q�q�?             (@       �       �                   �<@      �?              @        ������������������������       �                     �?        �       �                 X�,@@և���X�?             @       �       �                 �|Y=@      �?             @        ������������������������       �                     �?        �       �                 `fF<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 03k:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    R@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��|�5��?            �G@       �       �                 `ށK@���y4F�?             C@       �       �                    �?�IєX�?             1@       �       �                    �?$�q-�?
             *@        ������������������������       �                     @        �       �                 �|�<@ףp=
�?             $@        �       �                 `f�D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 X��@@�q�q�?
             5@        ������������������������       �                     $@        �       �                   �H@���|���?             &@       �       �                   @G@      �?              @        �       �                   �D@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�q�q�?             "@       �       �                    �?�q�q�?             @       �       �                    �?      �?             @       �       �                 03/O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    /@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �                       �T�I@įDg50�?=            @Y@       �       �                    0@NKF����?7            @V@        �       �                   �/@���Q��?             4@       �       �                   �-@�t����?             1@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �5@d}h���?	             ,@        ������������������������       �                     �?        �       �                    �?8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��d2@�LQ�1	�?+            @Q@        ������������������������       �                     (@        �       �                    �?�S����?%            �L@        �       �                    �?      �?              @       �       �                 м;4@�q�q�?             @        �       �                   �2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                          @�q��/��?            �H@       �                       ��T?@��E�B��?            �G@                                 @l��\��?             A@        ������������������������       �                      @                                 �?      �?             @@       ������������������������       �                     8@                                  @      �?              @        ������������������������       �                     �?                                 �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        	                         �?�θ�?             *@       
                        �C@�C��2(�?             &@                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @                                  @�q�q�?             (@        ������������������������       �                     @                              p�O@�<ݚ�?             "@                                >@      �?              @                                ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������N���I5�?d�~`l��?1�0��?�y��y��?���(0��?���g��?��,d!�?8��Moz�?��y��y�?�a�a�?�m۶m۶?I�$I�$�?"5�x+��?��sHM0�?      �?      �?      �?      �?      �?                      �?              �?l�l��??�>��?              �?�������?�������?              �?�������?333333�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?)\���(�?�Q����?��,d!�?8��Moz�?t�E]t�?��.���?              �?�������?ZZZZZZ�?      �?      �?              �?�������?�������?      �?                      �?      �?        ��+��+�?����?��y��y�?�a�a�?�������?�������?      �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?              �?�$I�$I�?۶m۶m�?333333�?�������?              �?�+Q��?ە�]���?�{a���?��=���?UUUUUU�?UUUUUU�?ffffff�?333333�?9��8���?�q�q�?              �?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?              �?      �?              �?        ��8��8�?�q�q�?      �?        ]t�E�?F]t�E�?              �?      �?                      �?�A^%���?���j�1�?�.���?ݘ��V��?              �?����=	�?�gPE!l�?&�X�%�?O贁N�?۶m۶m�?�$I�$I�?      �?        333333�?333333�?�������?�?              �?n۶m۶�?�$I�$I�?      �?              �?      �?      �?              �?      �?�������?�������?              �?      �?        ����?���?      �?        ���k(�?(�����?*�Y7�"�?к����?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        .���r��?�F��h4�?��:��?XG��).�?۶m۶m�?�$I�$I�?      �?                      �?ܯK*��?���ϱ?%I�$I��?۶m۶m�?      �?        �<%�S��?�־a�?�������?�?�؉�؉�?;�;��?;�;��?;�;��?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?      �?              �?        6��P^C�?(������?              �?<<<<<<�?�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ��N��?'u_[�?�/����?�}A_Ч?      �?        ӛ���7�?d!Y�B�?      �?        �������?UUUUUU�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?        �������?�������?              �?      �?        0&q��?ӟ���?ffffff�?333333�?e�M6�d�?N6�d�M�?۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?�$I�$I�?۶m۶m�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?�������?      �?                      �?br1���?x6�;��?6��P^C�?(������?�?�?�؉�؉�?;�;��?      �?        �������?�������?      �?      �?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?        F]t�E�?]t�E]�?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        B���be�?�F�tj�?��g<��?�9�as�?333333�?�������?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?I�$I�$�?۶m۶m�?              �?;�;��?;�;��?      �?                      �?              �?��Moz��?Y�B��?      �?        (������?^Cy�5�?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        /����?և���X�?�l�w6��?AL� &W�?------�?�������?              �?      �?      �?      �?              �?      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?        ى�؉��?�؉�؉�?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?                      �?      �?        �������?�������?      �?        �q�q�?9��8���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ?{�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM#hjh))��}�(h,h/h0M#��h2h3h4hph<�h=Kub������       �                 `�X.@>AU`�z�?�           8�@               ?                    �?Z���,<�?�            v@               8                 P�>,@t�����?7             U@              3                    �?����?2            @S@                                 �5@��M���?,             Q@                                   �?$�q-�?	             *@        ������������������������       �                     @                                   �?      �?              @       	                          �3@r�q��?             @       
                        P��@      �?             @        ������������������������       �                      @                                ��!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                   �?��N`.�?#            �K@                                �|Y:@z�G�z�?             4@        ������������������������       �                     @                                   �?������?             1@        ������������������������       �                     �?                                ���@      �?             0@        ������������������������       �                     @                                ���@$�q-�?
             *@        ������������������������       �                      @                                   �?�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?               &                     @���Q��?            �A@                               `f�)@�r����?             .@        ������������������������       �                     @                !                    ;@      �?              @        ������������������������       �                     �?        "       #                   �B@؇���X�?             @       ������������������������       �                     @        $       %                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        '       0                 �|�=@���Q��?
             4@       (       +                    8@������?             .@        )       *                   �6@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ,       -                 �&B@�����H�?             "@        ������������������������       �                     @        .       /                    ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        1       2                 ��n @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        4       7                   �!@�q�q�?             "@        5       6                    6@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        9       :                    �?؇���X�?             @        ������������������������       �                     @        ;       >                 pF�,@      �?             @       <       =                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        @       �                    �?$Z�?�            �p@       A       R                    �?ĴF���?�            �n@        B       I                 �|Y=@lGts��?            �K@        C       H                 �Y�@և���X�?             @       D       E                    5@z�G�z�?             @        ������������������������       �                      @        F       G                   @9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        J       K                    �?      �?             H@       ������������������������       �                     9@        L       Q                 X�I@�LQ�1	�?             7@       M       N                  s�@��2(&�?             6@        ������������������������       �                     @        O       P                 ��(@r�q��?             2@       ������������������������       �@�0�!��?             1@        ������������������������       �                     �?        ������������������������       �                     �?        S       �                    �?��Y���?~            �g@       T       �                   @E@�>����?|            �g@       U       d                 �?�@ĴF���?m            �d@        V       W                   �7@ ���J��?4            �S@        ������������������������       �                     >@        X       c                 �?$@ �q�q�?#             H@        Y       Z                 �&b@�C��2(�?             6@        ������������������������       �                     (@        [       \                   �8@z�G�z�?             $@        ������������������������       �                     �?        ]       ^                 �|�;@�����H�?             "@        ������������������������       �                     @        _       b                 �|Y?@r�q��?             @       `       a                 pf�@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     :@        e       l                 @3�@(L���?9            �U@        f       g                    :@      �?             @        ������������������������       �                     �?        h       i                   �?@���Q��?             @        ������������������������       �                      @        j       k                   �A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        m       �                    D@���(\��?4             T@       n       �                    &@���Lͩ�?1            �R@       o       �                 ���"@      �?%             L@       p       s                   �2@��-�=��?            �C@        q       r                 ��Y @����X�?             @        ������������������������       �                      @        ������������������������       �                     @        t       u                 ��) @      �?             @@       ������������������������       �                     5@        v       w                 ��y @"pc�
�?             &@        ������������������������       �                     �?        x                        @3"@ףp=
�?             $@       y       z                 pf!@z�G�z�?             @        ������������������������       �                     �?        {       ~                 �|Y<@      �?             @        |       }                    8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    $@@�0�!��?             1@       �       �                   �<@z�G�z�?             $@       ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    5@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     3@        �       �                     @���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     9@        �       �                   @7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    -@��<b���?             7@        ������������������������       �                     @        ������������������������       �                     2@        �       �                     @���$���?�            `v@       �       �                   �M@�4��?�            @p@       �       �                    �?~����?�            `n@       �       �                    @��<b�ƥ?T            @a@        �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    6@���%yU�?R            �`@        �       �                   @4@r�q��?             @       ������������������������       �                     @        �       �                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?����}��?M            �_@        ������������������������       �                     �J@        �       �                   �E@`׀�:M�?-            �R@       ������������������������       �        #            �N@        �       �                    �?$�q-�?
             *@        �       �                   @G@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�q�q�?F            @Z@       �       �                    �?ι�~��?8            �U@        �       �                 p�w@�z�G��?             >@       �       �                 p"�X@      �?             <@       �       �                   �;@8����?             7@        �       �                    �?�q�q�?             @       �       �                 ��LK@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    B@      �?             4@       �       �                 ���=@؇���X�?             ,@        �       �                    �?���Q��?             @       �       �                 �ܵ<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?      �?             @       �       �                    H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    :@      �?&             L@        ������������������������       �                      @        �       �                   �<@�q�q�?"             H@        �       �                    �?r�q��?             @       �       �                 `fF:@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?d}h���?             E@       �       �                   �G@�<ݚ�?             ;@       �       �                   @@@��2(&�?             6@        ������������������������       �                     "@        �       �                     �?�θ�?             *@       �       �                 `f�;@�z�G��?             $@       �       �                 03k:@      �?             @        ������������������������       �                     �?        �       �                   �C@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `f�<@���Q��?             @       �       �                     �?�q�q�?             @       �       �                    J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                     �?z�G�z�?             .@       �       �                   �E@�q�q�?             "@       �       �                   �B@      �?             @        ������������������������       �                      @        �       �                  x#J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �7@p�ݯ��?             3@        ������������������������       �                     "@        �       �                 �̾w@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                  )?@�t����?             1@        �       �                    R@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        �                          �?~	~���?@            �X@        �       �                    �?X�<ݚ�?             ;@        �       �                 ��.@�q�q�?	             .@        �       �                    �?r�q��?             @        ������������������������       �                     �?        �       �                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                 ��.@�q�q�?	             (@        ������������������������       �                     @        �                          @�<ݚ�?             "@       �                        �|�;@���Q��?             @        ������������������������       �                     �?                               �v6@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 0@�ˡ�5��?.            �Q@                                �4@      �?             @        ������������������������       �                      @              	                pff/@      �?             @        ������������������������       �                      @        
                         �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              "                   @��ɉ�?*            @P@                             ��T?@@�r-��?(            �M@                                �?�ʈD��?            �E@        ������������������������       �                     4@                                 4@�㙢�c�?             7@        ������������������������       �                     $@                              �̌4@�	j*D�?
             *@                                �B@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                 �?     ��?             0@                                 @      �?              @                                 ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @              !                   @      �?              @                              ��p@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M#KK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?s� ����?6v}3Y��?�y��y��?�0�0�?�S{��?
qV~B��?�������?�?;�;��?�؉�؉�?              �?      �?      �?UUUUUU�?�������?      �?      �?              �?      �?      �?      �?                      �?              �?              �?� O	��?��oX���?�������?�������?              �?�?xxxxxx�?              �?      �?      �?      �?        ;�;��?�؉�؉�?              �?F]t�E�?]t�E�?              �?      �?        �������?333333�?�?�������?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?wwwwww�?�?      �?      �?      �?                      �?�q�q�?�q�q�?      �?              �?      �?              �?      �?        �������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        ۶m۶m�?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ɡ.K5��?��U��?E�JԮD�?ە�]�ڵ?�<%�S��?�־a�?�$I�$I�?۶m۶m�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?        ��Moz��?Y�B��?��.���?t�E]t�?      �?        �������?UUUUUU�?ZZZZZZ�?�������?      �?              �?        o��2�|�?�d�h��?�Kh/��?h/�����?E�JԮD�?ە�]�ڵ?��-��-�?�A�A�?      �?        �������?UUUUUU�?]t�E�?F]t�E�?      �?        �������?�������?              �?�q�q�?�q�q�?      �?        �������?UUUUUU�?�������?�������?      �?              �?      �?      �?              �?        ⎸#��?w�qG��?      �?      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?ffffff�?�����̼?�6�i�?�K~��?      �?      �?}˷|˷�?�A�A�?�m۶m��?�$I�$I�?              �?      �?              �?      �?      �?        /�袋.�?F]t�E�?              �?�������?�������?�������?�������?      �?              �?      �?      �?      �?      �?                      �?      �?              �?        ZZZZZZ�?�������?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?        333333�?�������?      �?      �?      �?              �?              �?      �?              �?      �?        ��,d!�?��Moz��?              �?      �?        I=W�l�?\@aT���?�Z��Z��?�R+�R+�?�lC@�9�?�I�_c�?d!Y�B�?��7��M�?�������?�������?              �?      �?        ���̎?M�3�τ�?UUUUUU�?�������?              �?      �?      �?      �?                      �?�@ �?����~��?              �?к����?��L��?              �?;�;��?�؉�؉�?UUUUUU�?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?�w�q�?G�w��?ffffff�?333333�?      �?      �?d!Y�B�?8��Moz�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?      �?۶m۶m�?�$I�$I�?333333�?�������?      �?      �?      �?                      �?      �?              �?              �?      �?      �?      �?              �?      �?                      �?      �?                      �?      �?      �?      �?        �������?�������?UUUUUU�?�������?�������?�������?      �?                      �?              �?I�$I�$�?۶m۶m�?9��8���?�q�q�?��.���?t�E]t�?      �?        ى�؉��?�؉�؉�?ffffff�?333333�?      �?      �?              �?333333�?�������?              �?      �?              �?              �?        �������?333333�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?�������?�������?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?                      �?      �?              �?        Cy�5��?^Cy�5�?              �?ffffff�?333333�?      �?                      �?<<<<<<�?�?333333�?�������?      �?                      �?      �?        �)x9/�?h�����?�q�q�?r�q��?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?        �������?�������?              �?      �?                      �?�������?�������?              �?9��8���?�q�q�?333333�?�������?              �?      �?      �?      �?                      �?      �?        �RO�o��?H���@��?      �?      �?              �?      �?      �?      �?              �?      �?              �?      �?        �����?�����?'u_�?��c+���?A_���?�}A_з?      �?        �7��Mo�?d!Y�B�?      �?        vb'vb'�?;�;��?�������?�������?              �?      �?              �?              �?      �?      �?      �?      �?      �?              �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��}whG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM)hjh))��}�(h,h/h0M)��h2h3h4hph<�h=Kub������       |                     @"��p�?�           8�@               #                   �<@��+��?�            `s@                                   �?~�X��?D            �Y@                                  �?�KM�]�?&            �L@        ������������������������       �                     :@               	                    @�n`���?             ?@                                ��1V@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        
                          �9@ȵHPS!�?             :@       ������������������������       �                     2@                                  �;@      �?              @                                ��m1@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                  �+@      �?             G@        ������������������������       �        
             ,@                                   �?     ��?             @@                                 �8@b�2�tk�?             2@        ������������������������       �                     @                                   �?d}h���?             ,@        ������������������������       �                      @                                  �;@      �?             (@                                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                `f�D@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               "                    �?؇���X�?             ,@                !                    5@      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        $       ]                  x#J@��~����?{            �i@       %       V                  �>@~�u���?S            �a@       &       U                   �R@�^���U�?C            �\@       '       T                   @>@      �?B             \@       (       S                   �M@���|���?A            �[@       )       6                   �?@���g�?<            �Y@        *       5                    �?�������?             A@       +       2                 �|�=@���!pc�?            �@@       ,       -                    �?��.k���?
             1@        ������������������������       �                     @        .       1                     �?      �?             (@        /       0                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        3       4                    �?      �?             0@        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     �?        7       R                    @��z4���?*            @Q@       8       C                    �?�ʻ����?)             Q@        9       B                    �? 7���B�?             ;@       :       A                   �*@ �q�q�?             8@        ;       <                   �'@$�q-�?             *@        ������������������������       �                     @        =       >                   �B@�����H�?             "@       ������������������������       �                     @        ?       @                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        D       E                 `f�)@������?            �D@        ������������������������       �                      @        F       Q                   @E@<���D�?            �@@        G       P                    �?����X�?	             ,@       H       K                     �?���|���?             &@        I       J                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        L       O                    �?      �?              @       M       N                    C@�q�q�?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             3@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        W       Z                    �? 	��p�?             =@       X       Y                     �?���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        [       \                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       k                   HR@     ��?(             P@        _       j                 ��LP@�n_Y�K�?	             *@       `       i                    �?z�G�z�?             $@       a       b                    �?�q�q�?             @        ������������������������       �                      @        c       d                    �?      �?             @        ������������������������       �                     �?        e       f                   �C@�q�q�?             @        ������������������������       �                     �?        g       h                 �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        l       m                    �?��x_F-�?            �I@       ������������������������       �                    �B@        n       o                 X�,@@����X�?
             ,@        ������������������������       �                     @        p       u                    �?���|���?             &@        q       r                    �?�q�q�?             @        ������������������������       �                     �?        s       t                   �B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        v       {                 ��^@      �?              @       w       z                    �?؇���X�?             @       x       y                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        }       ~                 03�@���h0�?�            y@        ������������������������       �                     7@               �                    �?����X�?�            �w@        �       �                    �?f�<�>��?B            �]@        �       �                 �&�)@      �?             D@       ������������������������       �                     8@        �       �                    @      �?             0@       �       �                    �?���Q��?             .@       �       �                 03�-@X�Cc�?             ,@       �       �                    �?���!pc�?             &@       �       �                   �-@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y=@�θ�?/            �S@        �       �                 ؼC1@� �	��?             9@       �       �                    �?������?
             1@       �       �                   �7@r�q��?             (@        ������������������������       �                     @        �       �                 �Y�@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �x"@���Q��?             @        ������������������������       �                     �?        �       �                    7@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���7@      �?              @        �       �                   �2@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���@�NW���?!            �J@        �       �                 ���@r�q��?             (@        ������������������������       �                     @        �       �                 �|�=@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        �       �                 �|Y?@������?            �D@       �       �                    �?�X�<ݺ?             B@       �       �                    �?��?^�k�?            �A@        ������������������������       �                     @        �       �                    �?(;L]n�?             >@       �       �                 ���@`2U0*��?             9@        ������������������������       �                     @        �       �                 ��(@P���Q�?	             4@       ������������������������       ��X�<ݺ?             2@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @�θ�?�            @p@        �       �                    �?@�0�!��?             1@        ������������������������       �                     @        �       �                 ���A@d}h���?             ,@       �       �                     @�8��8��?	             (@       ������������������������       �                     @        �       �                    @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?TWi&Ĥ�?�            `n@        �       �                 ���5@     ��?)             P@       �       �                    �?r�q��?             H@       �       �                 P�@�n_Y�K�?            �C@        �       �                   �7@�q�q�?             (@       �       �                 ���@      �?              @        ������������������������       �                      @        �       �                    �?r�q��?             @       �       �                    4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��L&@l��
I��?             ;@       �       �                   �9@�t����?	             1@       ������������������������       �                     (@        �       �                 @3�@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 @3�/@���Q��?             $@        ������������������������       �                     @        �       �                    �?z�G�z�?             @       �       �                 ��1@      �?             @       �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �#@�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                   �;@      �?             @        ������������������������       �                     �?        �       �                    >@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        �       �                    #@d��ϸ�?s            `f@        �       �                 03>@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       (                   �?�t����?p            @e@       �       '                   �?��}���?d            @c@       �       �                 �?�@��� ��?`            �b@        �       �                 �|Y=@�.ߴ#�?&            �N@       ������������������������       �                     A@        �       �                 �|�=@�����H�?             ;@       �       �                 pf�@�S����?             3@        ������������������������       �                      @        �       �                  sW@���!pc�?             &@        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       $                   �?
�GN��?:             V@       �       �                 @3�@�w>�
��?6            �T@        �       �                    :@      �?              @        ������������������������       �                     @        �       �                   �A@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        �                         �2@�J�4�?1            �R@        �                         �1@���Q��?             .@       �                         �0@���!pc�?             &@       �                        pFD!@�z�G��?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     �?                              ��Y @      �?             @        ������������������������       �                     @        ������������������������       �                     �?                              �T)D@ףp=
�?*             N@                             ��) @,�+�C�?&            �K@        ������������������������       �                     9@        	      
                0SE @�r����?             >@        ������������������������       �                     �?                              `�X#@ܷ��?��?             =@                             ���"@�LQ�1	�?             7@                             @Q!@      �?
             0@        ������������������������       �                     @                              @3�!@�C��2(�?             &@                             �|Y<@      �?              @                                 8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                �<@����X�?             @        ������������������������       �                     @                              �|Y=@      �?             @        ������������������������       �                     �?                              �|�=@�q�q�?             @        ������������������������       �                     �?                                �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               !                   ;@���Q��?             @        ������������������������       �                     �?        "      #                �|�>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        %      &                ��y'@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     0@        �*       h�h))��}�(h,h/h0M)KK��h2h3h4hVh<�h=Kub������������J54v��?l�����?=���?ra�q�?*9/���?kch����?(�����?�k(���?              �?�c�1��?�9�s��?333333�?�������?              �?      �?        �؉�؉�?��N��N�?              �?      �?      �?333333�?�������?              �?      �?                      �?      �?      �?      �?              �?      �?9��8���?�8��8��?      �?        ۶m۶m�?I�$I�$�?              �?      �?      �?UUUUUU�?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?j6��bP�?+�' :_�?���ϴ�? 2ܫ`��?c:��,��?:��,���?      �?      �?]t�E]�?F]t�E�?^�	���?C����?�������?�������?F]t�E�?t�E]t�?�������?�?              �?      �?      �?�������?333333�?              �?      �?              �?              �?      �?              �?      �?              �?        %~F���?̵s���?�������?<<<<<<�?h/�����?	�%����?UUUUUU�?�������?;�;��?�؉�؉�?              �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�|����?������?      �?        |���?|���?�m۶m��?�$I�$I�?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?              �?              �?                      �?      �?                      �?              �?������?�{a���?�.�袋�?F]t�E�?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?              �?     ��?ى�؉��?;�;��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        �?�������?              �?�m۶m��?�$I�$I�?      �?        ]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?UK��a�?Vi+��<�?      �?        �m۶m��?�$I�$I�?�"h8���?��/���?      �?      �?              �?      �?      �?333333�?�������?%I�$I��?�m۶m��?F]t�E�?t�E]t�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ى�؉��?�؉�؉�?)\���(�?�Q����?�?xxxxxx�?UUUUUU�?�������?              �?�$I�$I�?�m۶m��?      �?                      �?�������?333333�?      �?              �?      �?              �?      �?              �?      �?      �?      �?      �?                      �?      �?        萚`���?�x+�R�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?        p>�cp�?������?��8��8�?�q�q�?_�_��?�A�A�?      �?        �������?�?���Q��?{�G�z�?      �?        ffffff�?�������?��8��8�?�q�q�?      �?              �?                      �?      �?        ى�؉��?�؉�؉�?�������?ZZZZZZ�?              �?۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?        ��lC@��?w�M��:�?      �?      �?UUUUUU�?UUUUUU�?;�;��?ى�؉��?�������?�������?      �?      �?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?        Lh/����?h/�����?<<<<<<�?�?      �?        333333�?�������?              �?      �?        �������?333333�?              �?�������?�������?      �?      �?      �?      �?      �?                      �?      �?              �?        �q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �e㛡��?�ir�y)�?r�q��?�q�q�?              �?      �?        <<<<<<�?�?j`���?V~B����?��Ug��?7`��c.�?�K�`m�?XG��).�?      �?        �q�q�?�q�q�?(������?^Cy�5�?      �?        F]t�E�?t�E]t�?�������?333333�?      �?              �?        �E]t��?�袋.��?%����?��k���?      �?      �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?�z�G��?{�G�z�?333333�?�������?F]t�E�?t�E]t�?ffffff�?333333�?      �?      �?      �?              �?              �?      �?              �?      �?        �������?�������?�}��7��?��)A��?      �?        �������?�?              �?��=���?a���{�?��Moz��?Y�B��?      �?      �?      �?        ]t�E�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �m۶m��?�$I�$I�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        333333�?�������?              �?      �?      �?      �?                      �?�������?�������?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�,�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM#hjh))��}�(h,h/h0M#��h2h3h4hph<�h=Kub������       ^                    �?���$ӡ�?�           8�@                                   �?�6i����?�            �m@                                   @�m(�X�?8            @U@                               ��.@@4և���?7             U@                                   &@r�q��?             B@        ������������������������       �                     �?                                    @؇���X�?            �A@        ������������������������       �                      @        	                           �?�+$�jP�?             ;@        
                           �?�z�G��?             $@                                  �?r�q��?             @        ������������������������       �                     @                                �|Y6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?      �?             @        ������������������������       �                     �?                                �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                ���@�t����?             1@        ������������������������       �                     �?                                �|�9@      �?             0@        ������������������������       �                     @                                   �?ףp=
�?	             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     H@        ������������������������       �                     �?               W                 �D�H@���p9W�?f             c@              T                    �?Ɣ��Hr�?O            �]@               O                 0#
9@�O��i�?C            �Y@       !       D                    �?؀�:M�?2            �R@       "       C                 ���1@X�Emq�?$            �J@       #       ,                     @      �?"             H@        $       %                   �:@�z�G��?             4@        ������������������������       �                      @        &       +                    L@�<ݚ�?             2@       '       *                   �C@      �?             0@        (       )                   �B@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        -       <                    �?և���X�?             <@       .       ;                 `��!@�G�z��?             4@       /       0                 ���@     ��?             0@        ������������������������       �                     @        1       :                 `�X!@�eP*L��?	             &@       2       7                   �9@      �?              @       3       4                    5@z�G�z�?             @        ������������������������       �                      @        5       6                   �6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        8       9                 �|�;@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        =       >                 �!@      �?              @        ������������������������       �                      @        ?       @                 �|�;@      �?             @        ������������������������       �                      @        A       B                 ���.@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        E       F                    �?���N8�?             5@        ������������������������       �                     $@        G       N                 ��97@�eP*L��?             &@       H       I                     @؇���X�?             @        ������������������������       �                     @        J       M                    >@      �?             @       K       L                 P��%@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        P       Q                   @D@\-��p�?             =@       ������������������������       �                     4@        R       S                   @H@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        U       V                 ���0@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        X       Y                    �?г�wY;�?             A@       ������������������������       �                     <@        Z       ]                     @r�q��?             @        [       \                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        _       �                 `ff:@"��S�&�?           �}@       `       �                 `�X.@0��QQX�?�            �u@       a       b                    ,@8��8���?�             r@        ������������������������       �                     @        c       �                   @E@4_�����?�            �q@       d       �                    �?<��.���?�            �o@       e       f                     �?��I�?�             o@        ������������������������       �                     @        g       �                   @C@ i���t�?�            �n@       h       �                    �?�W�a=�?�            �l@       i       |                 �Y�@@݈g>h�?�            �l@        j       k                     @t/*�?            �G@        ������������������������       �                     @        l       w                   �8@��s����?             E@        m       r                    �?      �?             (@        n       o                 ���@      �?             @        ������������������������       �                      @        p       q                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        s       t                    7@      �?              @       ������������������������       �                     @        u       v                 �&b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        x       {                 �|�=@��S�ۿ?             >@       y       z                 ���@      �?             0@       ������������������������       �                     "@        ������������������������       �����X�?             @        ������������������������       �                     ,@        }       ~                  ��@�����?r            �f@        ������������������������       �                     3@               �                 �?$@|E+�	��?g            @d@        �       �                    �?���y4F�?             3@       �       �                 �|Y=@d}h���?
             ,@        ������������������������       �                     �?        �       �                    �?8�Z$���?	             *@       ������������������������       �"pc�
�?             &@        ������������������������       �                      @        �       �                 �|Y9@z�G�z�?             @       ������������������������       �                     @        ������������������������       �      �?              @        �       �                   �0@�'g�2�?X            �a@        ������������������������       ��q�q�?             @        �       �                     @ >�֕�?V            �a@        �       �                 ��,@HP�s��?             9@       �       �                 `fF)@�C��2(�?             6@       �       �                    &@@4և���?             ,@       �       �                   �5@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @@      �?              @        ������������������������       �                     @        �       �                   �A@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�=@P���Q�?C            �\@       �       �                 �?�@��V�I��?4            �W@        ������������������������       �                    �C@        �       �                    �?�1�`jg�?            �K@        ������������������������       �                     @        �       �                 @3�@0G���ջ?             J@        �       �                   �4@      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �9@ �q�q�?             H@        ������������������������       �                     ;@        �       �                   �;@�����?             5@        ������������������������       �                     �?        �       �                 pf� @P���Q�?             4@        �       �                 ��) @      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?؇���X�?             5@        ������������������������       �                     @        �       �                   �@@�0�!��?             1@        ������������������������       �                     �?        �       �                 ��)"@      �?             0@       �       �                   �?@��S�ۿ?             .@        �       �                   �>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             (@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �C@������?             .@        ������������������������       �      �?             @        �       �                     @�����H�?             "@        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     =@        �       �                    �?��mo*�?$            �M@        �       �                    /@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     �?D>�Q�?              J@        ������������������������       �                      @        �       �                    �?j�q����?             I@        �       �                   `3@؇���X�?             @        ������������������������       �                     @        �       �                 03�7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �̌4@&^�)b�?            �E@        �       �                     @j���� �?             1@        ������������������������       �                     @        �       �                 `f^4@����X�?
             ,@       �       �                    )@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �? ��WV�?             :@       ������������������������       �        
             4@        �       �                    ,@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �                          �?�j�'7m�?G            �_@       �       �                 03�I@@�&b
}�?0            �U@       �       �                    �?�F�j��?            �J@        �       �                 `f&;@�n_Y�K�?             *@        ������������������������       �                     @        �       �                   �A@      �?             $@       �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�=@z�G�z�?             @       �       �                 ��2>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 ��Y>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     �?�G�z��?             D@       �       �                   �B@��
ц��?            �C@       �       �                   �<@��.k���?             A@        ������������������������       �                     "@        �       �                 �|Y=@��H�}�?             9@        ������������������������       �                     @        �       �                  i?@8�A�0��?             6@       �       �                 `fF<@��.k���?
             1@       �       �                   �J@���!pc�?             &@       �       �                    H@      �?              @       �       �                 �|�?@����X�?             @        ������������������������       �                      @        �       �                   �C@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?                                   @�!���?             A@                                �?d��0u��?             >@                               �}S@z�G�z�?             .@        ������������������������       �                      @                               �	U@և���X�?             @        ������������������������       �                      @                                �5@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        	                         �?��S���?
             .@       
                        �E@�n_Y�K�?	             *@                             �w|c@      �?              @                               �B@����X�?             @                             `f�O@�q�q�?             @                                @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @              "                @�:x@R���Q�?             D@                                �?�L���?            �B@                                �4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                  @`Jj��?             ?@        ������������������������       �                     $@              !                   @�����?             5@                                 @�r����?
             .@        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M#KK��h2h3h4hVh<�h=Kub������������H�1�N�?oݟ�Kb�?T:�g *�?kq�w��?�?]]]]]]�?�$I�$I�?n۶m۶�?UUUUUU�?�������?      �?        �$I�$I�?۶m۶m�?              �?B{	�%��?/�����?333333�?ffffff�?UUUUUU�?�������?              �?      �?      �?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �?<<<<<<�?      �?              �?      �?              �?�������?�������?              �?      �?                      �?      �?        ������?������?#h8����?��c+���?��,��?�����?v�)�Y7�?E>�S��?�}�	��?5�x+��?      �?      �?333333�?ffffff�?      �?        �q�q�?9��8���?      �?      �?�$I�$I�?�m۶m��?              �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?      �?              �?]t�E�?t�E]t�?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?              �?      �?      �?      �?              �?      �?      �?                      �?      �?        ��y��y�?�a�a�?              �?]t�E�?t�E]t�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?      �?      �?                      �?              �?      �?        �{a���?a����?              �?�q�q�?r�q��?      �?                      �?�������?�?              �?      �?        �?�?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?�ґ=Q�?x��	��?�|�>��?�G*;�?�������?�������?              �?FI�8S,�?ӵ8f��?6��f���?M&��d2�?�������?&sp볹?      �?        /�����?����X�?�V���?vI�ø_�?�P^Cy�?Cy�5��?�;����?W�+���?      �?        z��y���?�a�a�?      �?      �?      �?      �?              �?      �?      �?              �?      �?              �?      �?      �?              �?      �?      �?                      �?�������?�?      �?      �?      �?        �m۶m��?�$I�$I�?      �?        ]��ҟ��?�jc�?      �?        ?,R�n�?�n���?6��P^C�?(������?I�$I�$�?۶m۶m�?              �?;�;��?;�;��?/�袋.�?F]t�E�?      �?        �������?�������?      �?              �?      �?$T�ik��?�^���?UUUUUU�?UUUUUU�?��+��+�?�A�A�?q=
ףp�?{�G�z�?]t�E�?F]t�E�?n۶m۶�?�$I�$I�?�q�q�?�q�q�?              �?      �?              �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?        �ø_�T�?��s���?<�����?AL� &W�?      �?        A��)A�?�־a�?      �?        vb'vb'�?�؉�؉�?      �?      �?      �?      �?      �?                      �?      �?        �������?UUUUUU�?      �?        =��<���?�a�a�?              �?ffffff�?�������?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?        ZZZZZZ�?�������?              �?      �?      �?�������?�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        wwwwww�?�?      �?      �?�q�q�?�q�q�?�������?�������?      �?              �?              �?        �<�"h�?W'u_�?�$I�$I�?�m۶m��?      �?                      �?b'vb'v�?vb'vb'�?      �?        =
ףp=�?
ףp=
�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���/��?�}A_��?�������?ZZZZZZ�?              �?�m۶m��?�$I�$I�?�������?�������?              �?      �?              �?      �?      �?                      �?O��N���?;�;��?      �?        �������?UUUUUU�?              �?      �?        �D"�H$�?�v��n��?�C��:��?)^ ���?��sHM�?:�&oe�?ى�؉��?;�;��?              �?      �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?�������?�������?�;�;�?�؉�؉�?�?�������?              �?{�G�z�?
ףp=
�?      �?        颋.���?/�袋.�?�?�������?F]t�E�?t�E]t�?      �?      �?�m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?      �?              �?      �?                      �?      �?              �?              �?        �������?�������?wwwwww�?DDDDDD�?�������?�������?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?�?�������?;�;��?ى�؉��?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?              �?                      �?              �?333333�?333333�?}���g�?L�Ϻ��?�������?UUUUUU�?              �?      �?        ���{��?�B!��?      �?        =��<���?�a�a�?�������?�?              �?      �?              �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�%\hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       �                    �?�,�٧��?�           8�@              �                  x#J@�U��F��?E           X�@              :                    �?���};��?           �{@                                `fV$@
�cՔ��?I            @^@                                   �?
j*D>�?              J@                                �|Y8@�C��2(�?             6@        ������������������������       �                     @                                ���@�����H�?             2@        	       
                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             ,@                                  �7@�q�q�?             >@                                  �?��.k���?
             1@                               pff@�q�q�?             (@                                  4@�����H�?             "@                                P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   4@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                �|�;@$�q-�?             *@                                  �9@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               9                    G@2L�����?)            @Q@              *                    �?     ��?&             P@                '                   �B@(N:!���?            �A@       !       "                    �?��S�ۿ?             >@        ������������������������       �                     @        #       &                   �9@�8��8��?             8@        $       %                   �6@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             2@        (       )                   �*@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        +       4                 03�1@д>��C�?             =@       ,       /                   �-@�t����?             1@        -       .                   �,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        0       1                 �|Y<@��S�ۿ?	             .@        ������������������������       �                     @        2       3                  S�-@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        5       6                    6@      �?	             (@        ������������������������       �                      @        7       8                   �E@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ;       �                    �?�Zl�i��?�            @t@       <       K                     �?���	���?�            r@        =       >                   �@@� ��1�?            �D@        ������������������������       �        
             .@        ?       @                 ��$:@�	j*D�?             :@        ������������������������       �                     @        A       B                   @E@D�n�3�?             3@        ������������������������       �                     @        C       J                    R@d}h���?	             ,@       D       I                 `f�;@8�Z$���?             *@       E       H                   �J@      �?              @       F       G                    H@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        L       M                 ���@x��A��?�             o@        ������������������������       �                     ;@        N       k                 �|Y=@�ͳ ���?�            �k@        O       P                 03�@fGk�T�?=            �W@        ������������������������       �                     @        Q       R                     @�A����?;             W@        ������������������������       �        
             *@        S       T                 ���@p#�����?1            �S@        ������������������������       �                     (@        U       f                   �<@� y���?)            �P@       V       W                 �?�@ܷ��?��?$             M@        ������������������������       �                     3@        X       e                 @�!@8�Z$���?            �C@       Y       d                   �:@�+e�X�?             9@       Z       c                   �3@�㙢�c�?             7@       [       `                   �2@������?	             .@       \       _                 ��Y @z�G�z�?             $@        ]       ^                    1@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        a       b                 0S5 @���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             ,@        g       h                    �?X�<ݚ�?             "@        ������������������������       �                     @        i       j                 ���"@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        l       {                   �@@4և���?R            �_@        m       t                 ��@�Ra����?             F@       n       s                 �|�=@г�wY;�?             A@       o       r                 �Y�@XB���?             =@        p       q                 ���@�����H�?             "@        ������������������������       �                     @        ������������������������       �z�G�z�?             @        ������������������������       �        
             4@        ������������������������       �                     @        u       v                    �?���Q��?             $@        ������������������������       �                      @        w       z                 �&B@      �?              @       x       y                 �|Y>@և���X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        |       }                 �|�=@������?5            �T@        ������������������������       �                     @@        ~       �                   �?@HP�s��?#             I@               �                     @����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �? �#�Ѵ�?            �E@        ������������������������       �                      @        �       �                 `fF)@ >�֕�?            �A@        ������������������������       �                     4@        �       �                   �*@�r����?             .@       �       �                   �F@      �?              @       �       �                   �A@���Q��?             @        ������������������������       �      �?              @        �       �                   �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��?^�k�?            �A@        �       �                     @�8��8��?             (@        ������������������������       �                     @        �       �                 �|Y<@؇���X�?             @        ������������������������       �                      @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     7@        �       �                 03?U@���B���?-            �S@        �       �                    �?">�֕�?            �A@        �       �                    �?�t����?
             1@       ������������������������       �                     &@        �       �                   �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     @      �?
             2@       �       �                    >@��S���?             .@        ������������������������       �                     @        �       �                 03�M@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �2@�ʈD��?            �E@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �H@��p\�?            �D@       �       �                 �|�=@�}�+r��?             C@        �       �                    �?r�q��?
             (@        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     :@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���t���?n            �g@       �       �                    �?���!pc�?A            �[@        �       �                 �|Y>@�?�P�a�?              N@       �       �                     @>A�F<�?             C@        ������������������������       �        	             3@        �       �                    @p�ݯ��?
             3@        ������������������������       �                      @        �       �                    �?���|���?             &@        ������������������������       �                      @        �       �                    �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     6@        �       �                 ��97@z�):���?!             I@        �       �                     @ףp=
�?             $@        ������������������������       �                     @        �       �                    �?r�q��?             @       �       �                    @�q�q�?             @       �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @�G�z��?             D@        �       �                 ���[@r�q��?             2@       ������������������������       �                     "@        �       �                    $@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    @��2(&�?             6@       ������������������������       �                     *@        �       �                    @�q�q�?             "@        �       �                 ��T?@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    :@����?-            �S@        �       �                    �?r�q��?             8@       �       �                    �?�\��N��?             3@        ������������������������       �                     @        �       �                    �?     ��?             0@       �       �                    #@      �?
             ,@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     @PN��T'�?             K@       �       �                     �?x�����?            �C@       �       �                   �4@�+e�X�?             9@        ������������������������       �                     @        �       �                    �?�����?	             5@       �       �                 �̾w@�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?؇���X�?             ,@       �       �                    0@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             .@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������&��jq�?:�g *�?�Zؒ��?��KO��?y1��%��?����?"pc�
�?�GN�z�?;�;��?b'vb'v�?F]t�E�?]t�E�?              �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?�?�������?UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?        �������?�������?              �?      �?        �؉�؉�?;�;��?�������?UUUUUU�?      �?                      �?      �?        �Q�g���?�k�ځ�?      �?     ��?�A�A�?|�W|�W�?�?�������?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?333333�?      �?                      �?|a���?a���{�?�?<<<<<<�?      �?      �?              �?      �?        �?�������?              �?�������?�������?      �?                      �?      �?      �?      �?        �������?�������?              �?      �?              �?        �"e����?�����H�?d��E��?:߄*�u�?������?������?      �?        vb'vb'�?;�;��?      �?        l(�����?(������?              �?I�$I�$�?۶m۶m�?;�;��?;�;��?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?!�B�?���{ｷ?      �?        ]p�\p��?}�}��?��c�H�?�-q����?              �?C���,�?�Mozӛ�?      �?        7a~W��?�#{���?      �?        z�rv��?~5&��?��=���?a���{�?      �?        ;�;��?;�;��?R���Q�?���Q��?�7��Mo�?d!Y�B�?wwwwww�?�?�������?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?              �?                      �?      �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?                      �?n۶m۶�?�$I�$I�?]t�E]�?]t�E�?�?�?GX�i���?�{a���?�q�q�?�q�q�?      �?        �������?�������?      �?              �?        333333�?�������?      �?              �?      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?p>�cp�?������?      �?        q=
ףp�?{�G�z�?�m۶m��?�$I�$I�?      �?                      �?�/����?�}A_Ч?      �?        ��+��+�?�A�A�?      �?        �������?�?      �?      �?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?        _�_��?�A�A�?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?      �?        ى�؉��?��؉���?�A�A�?_�_��?�?<<<<<<�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�?�������?      �?        F]t�E�?]t�E]�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�}A_з?A_���?      �?      �?              �?      �?        ��+Q��?�]�ڕ��?(�����?�5��P�?UUUUUU�?�������?�������?333333�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?���\AL�?���Q���?t�E]t�?F]t�E�?�����ݽ?DDDDDD�?Cy�5��?������?              �?Cy�5��?^Cy�5�?              �?]t�E]�?F]t�E�?              �?9��8���?�q�q�?              �?      �?                      �?q=
ףp�?H�z�G�?�������?�������?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?�������?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?��.���?t�E]t�?      �?        UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?      �?        H�4H�4�?��-��-�?UUUUUU�?UUUUUU�?�5��P�?y�5���?              �?      �?      �?      �?      �?              �?      �?              �?        �������?�������?      �?                      �?&���^B�?h/�����?��o��o�?�A�A�?R���Q�?���Q��?              �?=��<���?�a�a�?�������?�?      �?                      �?      �?        ۶m۶m�?�$I�$I�?9��8���?�q�q�?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ2�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                  x#J@"��p�?�           8�@              [                    �?��n:���?w           ��@                                   �?P�|

��?z             h@                                �?�-@���5��?            �L@                               P�>,@     ��?             @@                               �|Y:@ ��WV�?             :@        ������������������������       �                     "@                                ���@�IєX�?
             1@        	       
                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     @        ������������������������       �                     9@               &                  �#@�>z���?[             a@               %                    �?���Q��?             4@                               ���@p�ݯ��?             3@        ������������������������       �                     @               $                    �?      �?             0@              #                    A@�q�q�?             (@              "                 �|Y>@X�<ݚ�?	             "@              !                    ;@      �?              @                                03�!@      �?             @                               �&B@���Q��?             @                                  �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                P�@�q�q�?             @        ������������������������       �                     �?                                  �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        '       Z                    @�������?K             ]@       (       E                   �?@p9W��S�?I            �\@       )       >                    �?2lK����?4            @T@       *       1                    7@d��0u��?&             N@        +       0                    �?(;L]n�?             >@        ,       -                     @�8��8��?             (@       ������������������������       �                     $@        .       /                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        2       =                 039@���Q��?             >@       3       <                 ��Y1@      �?             8@       4       ;                 �|�<@�t����?
             1@       5       :                 `f�,@�n_Y�K�?             *@       6       9                    �?X�<ݚ�?             "@       7       8                   �9@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ?       @                     @����X�?             5@        ������������������������       �                     @        A       D                    @      �?             0@        B       C                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             ,@        F       U                     @6YE�t�?            �@@       G       T                    L@ܷ��?��?             =@       H       M                   �*@@4և���?             <@        I       J                    B@؇���X�?             @        ������������������������       �                     @        K       L                    F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        N       O                  ��9@���N8�?             5@       ������������������������       �                     ,@        P       S                    :@؇���X�?             @        Q       R                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        V       Y                    �?      �?             @       W       X                 `f�/@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        \       a                    @p?ܘ�j�?�            y@        ]       `                   �C@և���X�?             5@       ^       _                    @z�G�z�?	             .@       ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     @        b       c                 03�@\�����?�            �w@        ������������������������       �                    �B@        d       �                     @d���X��?�            pu@        e       �                   @R@�C��2(�?L            @^@       f       �                    �?�8��8��?K             ^@       g       �                   �J@W�!?�?>            �X@       h       �                   �H@,���i�?3            �T@       i       �                   �>@�s�c���?/            @S@       j       q                    �?�? Da�?&            �O@        k       p                    �?      �?              @       l       o                 �|�=@؇���X�?             @        m       n                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        r       �                 `f�<@X�;�^o�?!            �K@       s       �                    �?0��_��?             �J@       t                          �@@`�H�/��?            �I@       u       ~                 `fv3@�FVQ&�?            �@@       v       y                    5@�����?             5@        w       x                   �2@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        z       {                 �|�<@�IєX�?             1@       ������������������������       �                     "@        |       }                 �|�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                   @A@r�q��?             2@        ������������������������       �                      @        �       �                 03K3@      �?
             0@        �       �                   �'@r�q��?             @        ������������������������       �                     �?        �       �                   @D@z�G�z�?             @        ������������������������       �                      @        �       �                   �F@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             ,@        �       �                     �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                     5@        ������������������������       �                     �?        �       �                    @`�t�D7�?�            �k@       �       �                    �?�)j9�v�?�            `j@        �       �                   �7@����X�?            �A@        �       �                    �?؇���X�?             @       �       �                 xF*@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���@؇���X�?             <@        ������������������������       �                      @        �       �                 �|�=@z�G�z�?	             4@       �       �                   �<@�q�q�?             (@        ������������������������       �                     @        �       �                   @@      �?              @        ������������������������       �                      @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?h�V���?v             f@        �       �                   `3@H%u��?             9@       �       �                 �|Y=@P���Q�?             4@        �       �                    ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     1@        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?tX�}}��?f            �b@       �       �                    �?�\�)G�?X            �`@       �       �                 P�N@pJQg���?W            �`@        �       �                 �|�<@Pa�	�?            �@@       ������������������������       �                     8@        �       �                 ��@�����H�?	             "@       ������������������������       �                     @        �       �                 �|Y>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �Yu@H%u��??             Y@        �       �                    >@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�=@�ɮ����?;            �V@       �       �                 ���"@�g�y��?*             O@       �       �                   �3@`Ql�R�?            �G@        �       �                   �2@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     E@        �       �                 `�X#@��S�ۿ?             .@        �       �                   �<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �?@>���Rp�?             =@        �       �                 �?�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 @3�@�LQ�1	�?             7@        �       �                   @C@      �?             (@       ������������������������       �                     @        �       �                 �?�@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                      @        �       �                    )@      �?             0@        ������������������������       �                     �?        �       �                 03S&@��S�ۿ?             .@        �       �                    �?z�G�z�?             @       �       �                    �?�q�q�?             @       �       �                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             $@        ������������������������       �                     &@        �       �                    �?��Sݭg�?M            @]@       �       �                     @����Q8�?0            �Q@       ������������������������       �        -            �P@        ������������������������       �                     @        �       �                    2@\X��t�?             G@        ������������������������       �                     @        �       �                    �?�ՙ/�?             E@        �       �                   �7@      �?
             0@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �                            �?
j*D>�?             :@       �       �                   �L@�X����?             6@       �       �                    6@      �?             4@        ������������������������       �                     �?        �       �                    �?���y4F�?             3@       �       �                 p"�X@      �?
             0@       �       �                    �?z�G�z�?	             .@        ������������������������       �                     @        �       �                    A@�z�G��?             $@        ������������������������       �                     @        �       �                 `�iJ@      �?             @        ������������������������       �                      @        �       �                 03�U@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������J54v��?l�����?R�Ω��?\��c�x�?n����?I	9��?��Gp�?�}��?      �?      �?;�;��?O��N���?              �?�?�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�?�������?333333�?�������?^Cy�5�?Cy�5��?              �?      �?      �?UUUUUU�?UUUUUU�?r�q��?�q�q�?      �?      �?      �?      �?�������?333333�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?                      �?      �?              �?                      �?,�4�rO�?j��FX�?l(�����?�k(����?�<ݚ�?��a�2��?�������?�?�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?�������?333333�?      �?      �?�������?�������?ى�؉��?;�;��?r�q��?�q�q�?۶m۶m�?�$I�$I�?      �?                      �?      �?                      �?              �?      �?                      �?�m۶m��?�$I�$I�?              �?      �?      �?      �?      �?      �?                      �?      �?        e�M6�d�?'�l��&�?a���{�?��=���?�$I�$I�?n۶m۶�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?�a�a�?��y��y�?              �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �1����?�8�Q�G�?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?        tK��=��?a�+F�?      �?        �=�P�\�?k&{��?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?�v���?1ogH�۹?�����?8��18�?�����?�cj`?�������?AA�?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?        �־a��?J��yJ�?"5�x+��?�V�9�&�?�������?�?>����?|���?=��<���?�a�a�?      �?      �?      �?                      �?�?�?      �?              �?      �?              �?      �?              �?        �������?UUUUUU�?              �?      �?      �?�������?UUUUUU�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?              �?                      �?      �?        333333�?�������?              �?      �?              �?              �?                      �?l��W���?Nq��$�?hn�����?_Fb5\��?�m۶m��?�$I�$I�?�$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �袋.��?/�袋.�?)\���(�?���Q��?ffffff�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        333333�?�������?      �?                      �?�Hs�9��?˸e�2n�?�Ε$��?n�Q�ߦ�?���7G��?\�qA��?|���?|���?      �?        �q�q�?�q�q�?      �?              �?      �?              �?      �?        )\���(�?���Q��?UUUUUU�?UUUUUU�?      �?                      �?]��\���?�Q�Q�?��{���?�B!��?}g���Q�?W�+�ɕ?�������?�������?      �?                      �?      �?        �������?�?�������?�������?      �?                      �?      �?        �i��F�?GX�i���?UUUUUU�?UUUUUU�?      �?                      �?��Moz��?Y�B��?      �?      �?      �?        �������?333333�?      �?                      �?      �?              �?              �?      �?              �?�������?�?�������?�������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?              �?              �?        �i�i�?�|˷|��?��Vج?O�o�z2�?              �?      �?        !Y�B�?��Moz��?              �?�<��<��?�a�a�?      �?      �?      �?      �?      �?                      �?      �?        ;�;��?b'vb'v�?]t�E]�?�E]t��?      �?      �?      �?        (������?6��P^C�?      �?      �?�������?�������?              �?333333�?ffffff�?              �?      �?      �?              �?      �?      �?      �?                      �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��(.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       Z                     @e�L��?�           8�@               U                    �?����o��?�            Pr@              0                     �?L8���?�             j@              #                    �?��7Y��?J            �[@                                  ;@�):u��?1            @S@        ������������������������       �                      @                                   �?
;&����?,            @Q@                                �D@J@`2U0*��?             9@        	       
                 ���;@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             4@                                   �?�������?             F@                                  @@@�C��2(�?             &@        ������������������������       �                     @                                  �A@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @               "                   �B@r٣����?            �@@                                 �<@�LQ�1	�?             7@        ������������������������       �                      @               !                    R@����X�?             5@                               �|�?@���y4F�?             3@                                  @>@�C��2(�?             &@       ������������������������       �                     @                                  �>@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                `fF:@      �?              @        ������������������������       �                     @                                   @M@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        $       %                    �?�t����?             A@        ������������������������       �                     2@        &       /                    �?      �?             0@       '       *                    �?�q�q�?             .@        (       )                   �5@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        +       .                    D@ףp=
�?             $@        ,       -                   @A@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        1       B                    �?�Y �K�?F            @X@        2       3                    �?b�h�d.�?            �A@        ������������������������       �                     @        4       ?                    �?�n`���?             ?@       5       :                   �B@H%u��?             9@       6       9                    :@�X�<ݺ?             2@        7       8                   �6@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             ,@        ;       <                   �'@����X�?             @        ������������������������       �                     �?        =       >                    D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        @       A                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     @        C       T                    ,@Hn�.P��?-             O@       D       S                    �?�˹�m��?             C@       E       R                   �A@�L���?            �B@       F       G                    @ �Cc}�?             <@        ������������������������       �                     @        H       M                   �(@      �?             8@        I       L                    &@�C��2(�?             &@       J       K                   �7@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        N       O                 �|�<@8�Z$���?
             *@       ������������������������       �                     $@        P       Q                 �|�?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     8@        V       W                    �?�c�x��?6            @U@       ������������������������       �        #             L@        X       Y                    4@>���Rp�?             =@        ������������������������       �                     @        ������������������������       �                     6@        [       �                    �?v����?�             z@        \       u                    �? ��X��?G            �]@        ]       t                    �?��x_F-�?            �I@       ^       k                    �?��[�p�?            �G@       _       d                    �? >�֕�?            �A@        `       a                    �?r�q��?             @        ������������������������       �                     �?        b       c                 �|Y6@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        e       j                    �?XB���?             =@       f       g                 �|Y8@`2U0*��?             9@        ������������������������       �                     @        h       i                 ���@���N8�?             5@        ������������������������       �                     �?        ������������������������       �        
             4@        ������������������������       �                     @        l       s                    �?�q�q�?             (@       m       r                  S�2@      �?              @       n       o                    3@�q�q�?             @        ������������������������       �                      @        p       q                 �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        v                        03s@h��Q(�?+            �P@       w       ~                    �?�7��?            �C@       x       }                 ���@���}<S�?             7@       y       z                 03S@8�Z$���?             *@        ������������������������       �                      @        {       |                   �7@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     $@        ������������������������       �                     0@        �       �                 ��.@և���X�?             <@        �       �                    �?�θ�?             *@       �       �                    3@և���X�?             @        ������������������������       �                     @        �       �                 �|Y=@      �?             @        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    /@�r����?
             .@        ������������������������       �                     @        �       �                 �|�8@�<ݚ�?             "@        ������������������������       �                     �?        �       �                    �?      �?              @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @���I��?�            �r@        �       �                    @�<ݚ�?
             2@       ������������������������       �                     $@        �       �                 ��T?@      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        �       �                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?Df/��?�            �q@       �       �                    �?� ��?�             o@       �       �                 ���@؇���X�?�             l@        ������������������������       �                     :@        �       �                 ���@n����W�?}            �h@        ������������������������       �                     �?        �       �                   �0@��(����?|            �h@        �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?     ��?z             h@        �       �                 �|�=@v�2t5�?            �D@       �       �                   �@���!pc�?            �@@        �       �                    �?�n_Y�K�?             *@       �       �                 �&B@�eP*L��?             &@       �       �                    8@      �?              @        �       �                 pf�@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|�<@P���Q�?             4@       ������������������������       �        	             .@        �       �                 pf&(@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�.(�i��?e            �b@       �       �                   �3@���۟�?^            `a@        �       �                 �?�@R���Q�?             4@       ������������������������       �                     (@        �       �                    2@      �?              @        ������������������������       �                     @        �       �                 �̌&@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 @Q!@�IєX�?S            �]@       �       �                 @3�@�ȉo(��?@            �V@       �       �                 �?�@��S�ۿ?,             N@       �       �                 �Yu@�&=�w��?&            �J@        �       �                 �|�<@�����?             5@       ������������������������       �        
             (@        �       �                 �&B@�<ݚ�?	             "@       �       �                 X�l@@      �?              @        �       �                 pf�@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @@        �       �                    :@����X�?             @        ������������������������       �                      @        �       �                   �?@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     ?@        �       �                   �;@ �Cc}�?             <@        �       �                    9@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                 �|�=@�X�<ݺ?             2@       ������������������������       �        	             ,@        �       �                 ��)"@      �?             @        ������������������������       �                      @        �       �                   @A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   �;@�+e�X�?             9@        �       �                    �?���|���?             &@        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                    @؇���X�?             @        �       �                 8�'@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?؇���X�?             ,@       �       �                 `fV6@z�G�z�?             $@        �       �                 `fv1@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    9@Pa�	�?            �@@        �       �                 ��L6@��S�ۿ?	             .@        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     2@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������v�S(��?��X��?���?wury�?;�;��?��؉���?\�9	ą�?�+c���?5�wL��?�'�Y�	�?              �?Y�B��?�Mozӛ�?{�G�z�?���Q��?�������?�������?              �?      �?                      �?t�E]t�?/�袋.�?]t�E�?F]t�E�?      �?        �������?UUUUUU�?              �?      �?        >���>�?|���?Nozӛ��?d!Y�B�?              �?�m۶m��?�$I�$I�?6��P^C�?(������?]t�E�?F]t�E�?      �?        �������?�������?              �?      �?              �?      �?      �?        �������?333333�?              �?      �?                      �?      �?        �������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?�������?�������?      �?      �?      �?                      �?      �?                      �?���
|q�?����?_�_��?;��:���?              �?�c�1��?�9�s��?���Q��?)\���(�?�q�q�?��8��8�?      �?      �?              �?      �?                      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?t�9�s�?�c�1ƨ?��P^Cy�?^Cy�5�?}���g�?L�Ϻ��?%I�$I��?۶m۶m�?      �?              �?      �?]t�E�?F]t�E�?۶m۶m�?�$I�$I�?      �?      �?      �?              �?        ;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?              �?        �������?�������?              �?�i��F�?GX�i���?              �?      �?        B�eh��?|�4�/��?qR���?[4���?�?�������?m�w6�;�?�
br1�?�A�A�?��+��+�?UUUUUU�?�������?              �?�������?�������?              �?      �?        �{a���?GX�i���?{�G�z�?���Q��?              �?�a�a�?��y��y�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?                      �?�Wc"=P�?z�rv��?��[��[�?�A�A�?ӛ���7�?d!Y�B�?;�;��?;�;��?      �?        /�袋.�?F]t�E�?              �?      �?              �?              �?        �$I�$I�?۶m۶m�?�؉�؉�?ى�؉��?۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?      �?                      �?      �?                      �?�������?�?      �?        9��8���?�q�q�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?Y�%�X�?�6�i��?�q�q�?9��8���?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?� &W��?G}g����?q����?<v5,���?۶m۶m�?�$I�$I�?      �?        )P�W
��?[�R�֯�?              �?��DO���?���b$�?�������?�������?              �?      �?             ��?      �?��+Q��?�ڕ�]��?F]t�E�?t�E]t�?ى�؉��?;�;��?]t�E�?t�E]t�?      �?      �?      �?      �?              �?      �?              �?                      �?              �?ffffff�?�������?      �?        �������?�������?      �?                      �?              �?���{��?��C�!��?��a����?����j�?333333�?333333�?      �?              �?      �?      �?              �?      �?              �?      �?        �?�?�~��?h�h��?�������?�?tHM0���?�x+�R�?=��<���?�a�a�?      �?        9��8���?�q�q�?      �?      �?      �?      �?      �?              �?      �?      �?                      �?      �?        �m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?      �?      �?        %I�$I��?۶m۶m�?�������?�������?      �?                      �?��8��8�?�q�q�?      �?              �?      �?      �?              �?      �?              �?      �?              �?        R���Q�?���Q��?]t�E]�?F]t�E�?              �?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?                      �?      �?              �?        |���?|���?�������?�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJx�+hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       `                    �?��ϙLq�?�           8�@               S                    @Rm�:Y�?�            `l@              J                 ��T?@����{@�?�            `i@              I                 0C�>@:-�.A�?Z            �`@              >                   @B@���!pc�?Y            �`@              =                 039@��Xk�?N             \@              <                   �>@     ��?E             X@                                  �?��X��?>             U@        	                          �-@z�G�z�?             D@        
                           �?�q�q�?             @        ������������������������       �                     @                                  �,@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?��hJ,�?             A@       ������������������������       �                     :@                                   �?      �?              @                                  @����X�?             @                               �|Y=@r�q��?             @                                03�-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?               3                    �?�eP*L��?!             F@                                    @������?             >@                                `f�)@�����H�?             "@       ������������������������       �                     @                                  �+@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        !       0                   �;@�q�q�?             5@       "       #                    @     ��?             0@        ������������������������       �                     @        $       +                 8�!@�θ�?	             *@       %       &                 ���@ףp=
�?             $@        ������������������������       �                     @        '       (                   �7@      �?             @        ������������������������       �                      @        )       *                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ,       -                   P&@�q�q�?             @        ������������������������       �                     �?        .       /                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       2                 �|�=@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        4       ;                    @؇���X�?             ,@       5       :                    �?$�q-�?
             *@       6       7                     @      �?              @        ������������������������       �                     �?        8       9                 �|Y;@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �        	             0@        ?       H                     @�G�z��?             4@       @       E                    �?     ��?	             0@       A       B                   �H@"pc�
�?             &@       ������������������������       �                     @        C       D                 03�3@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        F       G                   @F@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        K       R                    @��.N"Ҭ?.            @Q@       L       M                    �? ��ʻ��?-             Q@       ������������������������       �        &            �M@        N       O                 p"$X@�����H�?             "@        ������������������������       �                     @        P       Q                    $@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        T       _                    @      �?             8@       U       V                      @�z�G��?             4@        ������������������������       �                      @        W       Z                    @�<ݚ�?	             2@        X       Y                 ��T?@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        [       \                    @$�q-�?             *@       ������������������������       �                     "@        ]       ^                    ,@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        a       �                     �?�}�)ڳ�?0           @~@        b       �                 @�:x@v�C��?>            �X@       c       x                    �?���!���?<            �W@        d       s                    �?�!���?             A@       e       f                 ��";@z�G�z�?             9@        ������������������������       �                     �?        g       n                 03/O@r�q��?             8@       h       m                    �?��S�ۿ?
             .@       i       l                 ��2>@ףp=
�?             $@        j       k                 ���<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        o       p                    9@�q�q�?             "@        ������������������������       �                     �?        q       r                 p"�W@      �?              @        ������������������������       �                      @        ������������������������       �                     @        t       w                    �?�q�q�?             "@       u       v                 �U�X@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        y       z                 ��$:@���Q��?&             N@        ������������������������       �                     @        {       �                   �<@X�<ݚ�?"             K@        |       �                 `��P@"pc�
�?             &@       }       ~                 `ffC@����X�?             @        ������������������������       �                     @               �                    7@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �>@8�$�>�?            �E@        �       �                 03k:@�eP*L��?             6@        ������������������������       �                     @        �       �                    R@�\��N��?             3@       �       �                 �|Y=@      �?
             0@        ������������������������       �                      @        �       �                    K@և���X�?	             ,@       �       �                 `fF<@      �?             (@       �       �                 �|�?@�q�q�?             "@        ������������������������       �                     @        �       �                   �C@      �?             @        ������������������������       �                      @        �       �                    H@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?؇���X�?             5@       �       �                 03�U@�}�+r��?             3@       ������������������������       �                     0@        �       �                 X��@@�q�q�?             @        ������������������������       �                     �?        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?,�����?�            x@        �       �                     @p�v>��?             �G@        �       �                 `��.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 pF�#@������?            �D@       �       �                    �?H�V�e��?             A@       �       �                   �6@�'�`d�?            �@@        �       �                 ��y@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y=@�>����?             ;@        �       �                   @@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���@�nkK�?             7@        ������������������������       �                     &@        �       �                 �|Y?@�8��8��?             (@       �       �                   @@      �?              @       ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?����X�?             @       �       �                 03�-@r�q��?             @        �       �                   �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �                           �?PV�,��?�             u@       �       �                    )@0�v���?�            `p@        ������������������������       �                     @        �       �                    �?0_�n~f�?�            0p@       �       �                    �?     ��?�             p@        �       �                  ��@$�q-�?             :@        ������������������������       �                     "@        �       �                 �|Y=@�t����?             1@        ������������������������       �                      @        ������������������������       �        
             .@        �       �                     @���.�6�?�            �l@        �       �                    4@`'�J�?             �I@        �       �                   �2@�q�q�?             @        ������������������������       �                      @        �       �                   �'@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                    �F@        �       �                 �|Y=@FC��=�?k            `f@       �       �                   �:@ p�/��?:            @V@       �       �                   �9@p��%���?/            @Q@       �       �                 ���@     �?+             P@        �       �                 ���@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �3@���#�İ?&            �M@        �       �                   �2@���}<S�?             7@        ������������������������       �                     "@        �       �                 0S5 @؇���X�?             ,@       �       �                 �?�@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                     B@        �       �                 d�"@@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �       �                   @@@ףp=
�?1            �V@       �       �                 �?�@8�Z$���?             J@        �       �                 �|�=@���N8�?             5@       �       �                  sW@��S�ۿ?             .@       �       �                 pf�@      �?              @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                 @3�@��a�n`�?             ?@        �       �                   �?@      �?             $@        ������������������������       �                      @        ������������������������       �      �?              @        �       �                 ��) @�����?             5@        ������������������������       �                     $@        �       �                 �|�>@"pc�
�?             &@       �       �                 pf� @      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @C@P�Lt�<�?             C@        ������������������������       �        	             1@        �       �                   �C@���N8�?             5@        �       �                 ��	0@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �        	             1@        ������������������������       �                     @              
                   �?�S����?2             S@                              pf� @�FVQ&�?            �@@                                 7@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 6@h�����?             <@       ������������������������       �                     0@              	                03�7@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@                                 @>��C��?            �E@                                �;@     ��?             0@                                  @؇���X�?             @        ������������������������       �                     @                                  @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                              ��T?@�q�q�?             "@        ������������������������       �                     @                                  @      �?             @                             ��yE@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                              `f2@ 7���B�?             ;@                                  @�q�q�?             @        ������������������������       �                     �?                                �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������Ӭ����?�X�>��?�>c8Z�?��`����?igJ��8�?&f-б�?��~5&�?���@���?t�E]t�?F]t�E�?�m۶m��?�$I�$I�?      �?      �?%I�$I��?n۶m۶�?ffffff�?ffffff�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?KKKKKK�?              �?      �?      �?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?              �?]t�E�?t�E]t�?�?wwwwww�?�q�q�?�q�q�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?�؉�؉�?ى�؉��?�������?�������?              �?      �?      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?�������?      �?                      �?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?      �?                      �?              �?              �?�������?�������?      �?      �?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?      �?                      �?      �?              �?        ہ�v`��?�3J���?�?�������?              �?�q�q�?�q�q�?              �?�������?�������?      �?                      �?      �?              �?      �?ffffff�?333333�?              �?9��8���?�q�q�?�������?333333�?      �?                      �?�؉�؉�?;�;��?      �?              �?      �?      �?                      �?      �?        h���eP�?a���i��?gH���?1ogH���?�+���?�٨�l��?�������?�������?�������?�������?              �?�������?UUUUUU�?�������?�?�������?�������?�������?�������?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        333333�?�������?      �?        r�q��?�q�q�?F]t�E�?/�袋.�?�$I�$I�?�m۶m��?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?6eMYS��?�5eMYS�?]t�E�?t�E]t�?              �?y�5���?�5��P�?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?      �?      �?                      �?              �?      �?                      �?۶m۶m�?�$I�$I�?�5��P�?(�����?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?vN�07-�?M��{F��?ڨ�l�w�?L� &W�?UUUUUU�?UUUUUU�?              �?      �?        �v%jW��?��+Q��?iiiiii�?ZZZZZZ�?6�d�M6�?'�l��&�?UUUUUU�?�������?      �?                      �?�Kh/��?h/�����?      �?      �?      �?                      �?�Mozӛ�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?      �?      �?�������?�������?      �?              �?              �?        �$I�$I�?�m۶m��?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?        $��m��?ݾ�z�<�?�2����?�i��?              �?e޵M��?�Q:�Ͱ?     ��?      �?�؉�؉�?;�;��?      �?        <<<<<<�?�?              �?      �?        ���7���?Y�B��?�������?�?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        V,���?R�&���?�G?�я�?p�\��?�g��%�?ہ�v`��?     ��?      �?�������?�������?      �?                      �?��N��?'u_[�?ӛ���7�?d!Y�B�?      �?        ۶m۶m�?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?        �������?�������?      �?                      �?      �?        �������?�������?;�;��?;�;��?��y��y�?�a�a�?�������?�?      �?      �?      �?              �?      �?      �?              �?        �c�1��?�s�9��?      �?      �?              �?      �?      �?=��<���?�a�a�?      �?        /�袋.�?F]t�E�?      �?      �?              �?      �?              �?        ���k(�?(�����?      �?        ��y��y�?�a�a�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?              �?        (������?^Cy�5�?>����?|���?�������?�������?              �?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        $�;��?qG�w��?      �?      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?	�%����?h/�����?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJH�SshG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       `                    �?�3)0�F�?�           8�@               _                 ��R@     ��?�             p@              J                   @B@!��)��?~             i@              =                    @�MWl��?i            `e@              "                   �4@h������?\            �b@               !                   �3@��+7��?              G@                                  �?RB)��.�?            �E@              	                     @z�G�z�?             D@        ������������������������       �                     3@        
                        P��+@�ՙ/�?             5@                                  �?      �?	             (@                                  1@�q�q�?             "@        ������������������������       �                     @                                  �2@      �?             @                                  �?���Q��?             @                               ��!@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?X�<ݚ�?             "@                               03�-@z�G�z�?             @                                 �0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                    &@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        #       $                     @�̐d��?<            @Z@        ������������������������       �                    �I@        %       .                    �?����|e�?             K@        &       +                    �?��
ц��?             *@       '       *                 `�@1@և���X�?             @       (       )                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ,       -                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        /       8                    �?�p ��?            �D@       0       7                 �|�;@�#-���?            �A@        1       6                 pf(@      �?             (@       2       3                 P�@ףp=
�?             $@       ������������������������       �                     @        4       5                   �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     7@        9       :                    �?      �?             @        ������������������������       �                      @        ;       <                 @3s(@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        >       I                 �|Y?@�z�G��?             4@       ?       @                    @�d�����?             3@        ������������������������       �                     @        A       H                 �|Y7@�q�q�?             (@       B       C                    @����X�?             @        ������������������������       �                     �?        D       G                    *@r�q��?             @       E       F                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        K       X                 03;@*;L]n�?             >@       L       M                    �?      �?             4@        ������������������������       �                     �?        N       W                    �?���y4F�?             3@       O       V                     @      �?
             0@       P       U                    �?؇���X�?             ,@       Q       R                   �C@"pc�
�?             &@        ������������������������       �                     �?        S       T                    L@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        Y       ^                    @z�G�z�?             $@        Z       ]                    �?      �?             @       [       \                 83F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        !            �K@        a       l                    *@���w�?1           p|@        b       c                    @�q�q�?            �@@       ������������������������       �                     5@        d       e                    �?�8��8��?	             (@        ������������������������       �                     @        f       g                    �?؇���X�?             @        ������������������������       �                     @        h       i                    @�q�q�?             @        ������������������������       �                     �?        j       k                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        m       �                    @���V�?           `z@       n       �                    @"�q�?           @z@       o       �                    �?�$�S��?           �y@        p       �                     �?p�}�ޤ�?/            @R@        q       x                 �|Y<@     ��?             @@        r       w                  "&d@�θ�?             *@       s       v                   �8@r�q��?             (@       t       u                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        y       �                 tՌs@���y4F�?             3@       z                           �?r�q��?             2@       {       |                   �A@�θ�?             *@        ������������������������       �                     @        }       ~                   @J@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?,���i�?            �D@       �       �                   �5@$G$n��?            �B@        ������������������������       �                     �?        �       �                    �?�����H�?             B@       �       �                     @`Jj��?             ?@        ������������������������       �                      @        �       �                 �|Y=@���}<S�?             7@        �       �                   @@����X�?             @        ������������������������       �                     @        �       �                 ��Y&@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     0@        �       �                    �?���Q��?             @       �       �                     @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �R@��bH�e�?�            0u@       �       �                 ��D:@XY����?�             u@       �       �                    �?p��V	ַ?�            �q@       �       �                 ���@p�����?�            �p@        ������������������������       �        !             G@        �       �                    �? �o�b��?�            `k@        �       �                   `3@ȵHPS!�?             :@       �       �                 �|Y=@���}<S�?             7@        ������������������������       �                     �?        �       �                    �?���7�?             6@       �       �                 X��A@�X�<ݺ?             2@       �       �                 ��(@      �?	             0@       ������������������������       �$�q-�?             *@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 03�7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|Y=@�0p<���?�             h@       �       �                 ���$@T��,��?E            @Y@       �       �                   �3@@	tbA@�?/            @Q@        �       �                   �2@���N8�?             5@       ������������������������       �                     &@        �       �                 �?�@ףp=
�?             $@        ������������������������       �                     @        �       �                 0S5 @z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      H@        �       �                     @      �?             @@       �       �                    �?HP�s��?             9@       �       �                    &@�C��2(�?             6@        �       �                    5@      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     @        ������������������������       �                     @        �       �                   �C@���}<S�?=             W@       �       �                    �?H0sE�d�?0            �R@       �       �                     @ ���g=�?+            @Q@        �       �                 `fF)@@4և���?
             ,@        ������������������������       �                     @        �       �                 �|�=@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �@X�;�^o�?!            �K@        �       �                 �|�>@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                   @C@�:�]��?            �I@       �       �                 @3�@ �q�q�?             H@        �       �                    ?@      �?             0@       ������������������������       �                      @        �       �                 �?�@      �?              @       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                     5@        �       �                    �?      �?&             J@       �       �                 `f�;@�7����?"            �G@        �       �                   �J@�q�q�?	             (@       �       �                 03k:@�����H�?             "@        ������������������������       �                     �?        �       �                   @G@      �?              @       �       �                   �C@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                     �?؇���X�?            �A@       �       �                 03�M@6YE�t�?            �@@       �       �                 ��9L@�>4և��?             <@       �       �                   �<@PN��T'�?             ;@        �       �                 `f�D@      �?             @        ������������������������       �                     �?        �       �                    7@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �C@���}<S�?             7@        ������������������������       �                     $@        �       �                  i?@8�Z$���?             *@        �       �                   `H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?ףp=
�?             $@       ������������������������       �                     @        �       �                 �K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������Rl���?�[�'��?      �?     ��?��w����?�#�6���?�YLg1�?:��,���?��Tb*1�?��jg���?Y�B��?zӛ����?���)k��?S֔5eM�?�������?�������?              �?�a�a�?�<��<��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?333333�?�������?      �?      �?      �?                      �?              �?              �?              �?r�q��?�q�q�?�������?�������?      �?      �?              �?      �?              �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?         �����?��	��	�?              �?	�%����?����K�?�;�;�?�؉�؉�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?��+Q��?Q��+Q�?_�_�?�A�A�?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?ffffff�?333333�?Cy�5��?y�5���?      �?        �������?�������?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�������?""""""�?      �?      �?      �?        (������?6��P^C�?      �?      �?�$I�$I�?۶m۶m�?F]t�E�?/�袋.�?      �?        �������?�������?              �?      �?                      �?      �?                      �?�������?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?[�%[�%�?�6i�6i�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�<:�o�?�.~��?�Fk�Fk�?]ʥ\ʥ�?�R�yY�?<�o�14�?�z��ի�?�
*T��?      �?      �?�؉�؉�?ى�؉��?UUUUUU�?�������?�������?333333�?      �?                      �?              �?      �?        6��P^C�?(������?�������?UUUUUU�?ى�؉��?�؉�؉�?      �?              �?      �?              �?      �?              �?                      �?�����?8��18�?к����?���L�?              �?�q�q�?�q�q�?���{��?�B!��?      �?        ӛ���7�?d!Y�B�?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?              �?        333333�?�������?      �?      �?      �?                      �?      �?              �?        ����_[�?PR� %�?�%�q�?ц�s�?�ϴ5�n�?_���?<2l7O�?B�<���?      �?        E�}O��?�a�]�?��N��N�?�؉�؉�?ӛ���7�?d!Y�B�?              �?�.�袋�?F]t�E�?��8��8�?�q�q�?      �?      �?�؉�؉�?;�;��?      �?              �?              �?        UUUUUU�?UUUUUU�?              �?      �?        ��3-�?�O�l.�?�]?[��?�F�tj�?�%~F��?ہ�v`��?��y��y�?�a�a�?      �?        �������?�������?      �?        �������?�������?      �?      �?      �?              �?              �?      �?q=
ףp�?{�G�z�?]t�E�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?              �?              �?        ӛ���7�?d!Y�B�?��b�/��?O贁N�?��(�3J�?ہ�v`��?n۶m۶�?�$I�$I�?      �?        ]t�E�?F]t�E�?              �?      �?        �־a��?J��yJ�?      �?      �?UUUUUU�?UUUUUU�?              �?}}}}}}�?�?�������?UUUUUU�?      �?      �?      �?              �?      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?              �?      �?]AL� &�?G}g����?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?      �?      �?      �?      �?              �?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?'�l��&�?e�M6�d�?�$I�$I�?�m۶m��?&���^B�?h/�����?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?ӛ���7�?d!Y�B�?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?              �?      �?              �?      �?                      �?      �?              �?              �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�8�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM-hjh))��}�(h,h/h0M-��h2h3h4hph<�h=Kub������       j                 `f�$@�_%����?�           8�@               )                    �?��G���?�            0p@                                ���@l��
I��?%             K@                                ��Y@�8��8��?             8@        ������������������������       �                     @                                  @9@�KM�]�?
             3@        ������������������������       �                     �?               	                    �?�X�<ݺ?	             2@        ������������������������       �                      @        
                           �?      �?             0@                               ���@@4և���?             ,@        ������������������������       �                     @                                �|=@؇���X�?             @        ������������������������       �                     @                                �|�=@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @               (                 �|Y?@��S���?             >@                               @3�@��
ц��?             :@        ������������������������       �                     @                                   �?
;&����?             7@                                03@�����H�?	             "@                                  �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               '                    �?d}h���?             ,@                                �|Y=@8�Z$���?
             *@                                pfF@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        !       "                    �?ףp=
�?             $@        ������������������������       �                     �?        #       &                 ��(@�����H�?             "@       $       %                    �?؇���X�?             @       ������������������������       �r�q��?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        *       g                    �?�0]�I�?�            �i@       +       P                 �|�=@|g�&��?~            `i@       ,       ?                 �Yu@H%u��?]            �b@        -       .                 ���@��n�?+            �R@        ������������������������       �                     2@        /       0                 ���@P̏����?            �L@        ������������������������       �                      @        1       8                   �7@�rF���?            �K@       2       5                 P�N@�E��ӭ�?             B@       3       4                    �?�������?             >@        ������������������������       �                     @        ������������������������       �                     7@        6       7                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        9       :                    �?�KM�]�?             3@        ������������������������       �                     �?        ;       <                 �|�<@�X�<ݺ?             2@       ������������������������       �                     &@        =       >                 ��,@؇���X�?             @       ������������������������       �                     @        ������������������������       �      �?              @        @       C                   �0@Х-��ٹ?2            �R@        A       B                 pFD!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        D       M                    �?���(-�?0            @R@       E       L                 0SE @0�,���?,            �P@       F       G                   �2@�7��?            �C@        ������������������������       �                     �?        H       I                    �?P�Lt�<�?             C@        ������������������������       �                      @        J       K                 ��) @������?             B@       ������������������������       �                    �A@        ������������������������       �                     �?        ������������������������       �                     <@        N       O                   �4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        Q       V                    �?Ȩ�I��?!            �J@        R       U                  SE"@���Q��?             @       S       T                    C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        W       X                      @      �?             H@        ������������������������       �                     @        Y       f                   �C@������?            �F@       Z       e                   @C@ҳ�wY;�?             A@       [       d                 ��)"@�c�Α�?             =@       \       c                   @@@���B���?             :@       ]       ^                 �?�@     ��?	             0@        ������������������������       �                     @        _       b                 @3�@�eP*L��?             &@       `       a                   �?@����X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �z�G�z�?             @        ������������������������       �                     &@        h       i                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        k                         �R@n��Η��?!           @|@       l       �                    �?p� ��?�            �w@        m       �                     @j�$��?n            �d@       n       �                    L@` A�c̭?A             Y@       o       �                    �?`�E���??            @X@       p       �                    �?XB���?&             M@       q       v                   �9@`Ӹ����?            �F@        r       s                    �?�����H�?             "@        ������������������������       �                      @        t       u                   �6@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        w       x                     �?������?             B@        ������������������������       �                     @        y       z                    �?XB���?             =@        ������������������������       �                      @        {       |                   �B@ 7���B�?             ;@       ������������������������       �        
             1@        }       ~                   �'@ףp=
�?             $@        ������������������������       �                     @               �                   �,@r�q��?             @        �       �                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             *@        ������������������������       �                    �C@        �       �                   �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @�eP*L��?-            �P@        �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                 pf�0@؇���X�?             @        ������������������������       �                     @        �       �                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    7@      �?&             L@        �       �                    �?�X�<ݺ?             2@        �       �                 �&�)@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        �       �                   �C@�\��N��?             C@       �       �                  ��8@����e��?            �@@       �       �                    �?r�q��?             8@       �       �                    �?�㙢�c�?             7@       �       �                  S�-@@4և���?             ,@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �>@�q�q�?             "@       �       �                    �?���Q��?             @       �       �                 �|Y=@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                     �?�c�����?�            �j@        �       �                   �;@:PZ(8?�?0            @R@        �       �                    �?؇���X�?             @        ������������������������       �                     �?        �       �                    7@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �R@���!pc�?,            �P@       �       �                   �J@      �?+             P@       �       �                   �B@�q�q�?              H@       �       �                   �H@l��[B��?             =@       �       �                    �?�LQ�1	�?             7@        �       �                   @@@      �?              @        ������������������������       �                     @        �       �                    B@�q�q�?             @        ������������������������       �                     �?        �       �                 ��Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �F@���Q��?             .@       �       �                 �|�?@�eP*L��?
             &@       �       �                   @>@և���X�?             @        ������������������������       �                     @        �       �                   `@@      �?             @        ������������������������       �                      @        �       �                 �|�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    D@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                  x#J@�KM�]�?             3@       ������������������������       �                     $@        �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �                    >@�q�q�?             @        ������������������������       �                      @        �       �                 03�M@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                      @        �       �                     @(�}���?S            `a@       �       �                    %@� y���?*            �P@        ������������������������       �                     @        �       �                    �?85�}C�?&            �N@       �       �                 �|�=@�ݜ�?            �C@        �       �                    �?������?	             .@        ������������������������       �                     �?        �       �                 �|�<@����X�?             ,@       �       �                   �'@r�q��?             (@        �       �                    5@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �? �q�q�?             8@        ������������������������       �                     @        �       �                   @D@���N8�?             5@       ������������������������       �                     &@        �       �                    G@ףp=
�?             $@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     6@        �       �                    @<ݚ�?)             R@        �       �                    �?      �?
             2@       �       �                    �?��S���?             .@        ������������������������       �                     @        �       �                 ��|2@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                    @�q�q�?             @       �       �                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �                          ;@PN��T'�?             K@        �                          �3@      �?             4@       �       �                    �?�C��2(�?             &@        �       �                    '@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?X�<ݚ�?             "@        ������������������������       �                     @                                 7@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @              	                   �?l��\��?             A@                              `fv2@      �?             @       ������������������������       �                      @        ������������������������       �                      @        
                      �TE@(;L]n�?             >@       ������������������������       �                     ;@                                 �?�q�q�?             @                             �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?              ,                   �?���@��?0            �R@                             ���X@������?,             Q@                                 �?XB���?             =@       ������������������������       �                     5@                                �D@      �?              @        ������������������������       �                     @                                 �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                 �?�n_Y�K�?            �C@                             03c@�KM�]�?             3@                               "�b@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@               '                   �?��Q��?             4@       !      &                   �?�eP*L��?             &@       "      #                   �?r�q��?             @        ������������������������       �                     @        $      %                  �B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        (      )                ��f`@�<ݚ�?             "@       ������������������������       �                     @        *      +                ���i@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M-KK��h2h3h4hVh<�h=Kub������������z���� �?@Bx��?#�u�)��?v�)�Y7�?Lh/����?h/�����?UUUUUU�?UUUUUU�?      �?        �k(���?(�����?              �?��8��8�?�q�q�?      �?              �?      �?n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?      �?              �?        �?�������?�؉�؉�?�;�;�?              �?Y�B��?�Mozӛ�?�q�q�?�q�q�?UUUUUU�?�������?              �?      �?                      �?I�$I�$�?۶m۶m�?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?        �q�q�?�q�q�?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?              �?                      �?      �?        ٚ��I��?���Iٚ�?��v���?��%f-�?)\���(�?���Q��?:m���?�K~���?      �?        ?���#�?��Gp�?              �?yJ���?�־a��?�q�q�?r�q��?�������?�������?              �?      �?              �?      �?              �?      �?        �k(���?(�����?              �?��8��8�?�q�q�?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?K~��K�?O贁N�?      �?      �?              �?      �?        ��իW��?�P�B�
�?Ez�rv�?g��1��?��[��[�?�A�A�?              �?���k(�?(�����?      �?        �q�q�?�q�q�?      �?                      �?      �?        �������?UUUUUU�?              �?      �?        +�R��?�	�[���?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?        wwwwww�?�?�������?�������?5�rO#,�?�{a���?��؉���?ى�؉��?      �?      �?      �?        t�E]t�?]t�E�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?              �?                      �?�������?�������?      �?              �?      �?              �?      �?        d�:Fq�?�u��\��?�.6���?�䣓�N�?��ˊ��?�M�_{�?���Q��?
ףp=
�?����??��W�?�{a���?GX�i���?l�l��??�>��?�q�q�?�q�q�?              �?�$I�$I�?۶m۶m�?              �?      �?        �q�q�?�q�q�?              �?�{a���?GX�i���?              �?h/�����?	�%����?              �?�������?�������?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?UUUUUU�?UUUUUU�?      �?                      �?t�E]t�?]t�E�?�������?�������?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?��8��8�?�q�q�?      �?      �?              �?      �?              �?        �5��P�?y�5���?6�d�M6�?e�M6�d�?UUUUUU�?�������?d!Y�B�?�7��Mo�?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?      �?              �?        �V�9�&�?:�&oe�?�W�^�z�?�P�B�
�?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?      �?                      �?F]t�E�?t�E]t�?      �?      �?UUUUUU�?UUUUUU�?���=��?GX�i���?Nozӛ��?d!Y�B�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?333333�?�������?]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?              �?      �?      �?      �?                      �?�k(���?(�����?      �?        9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?U�wЍ�?�&!����?z�rv��?~5&��?              �?�}�K�`�?������?\��[���?�i�i�?wwwwww�?�?      �?        �m۶m��?�$I�$I�?�������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?                      �?�������?UUUUUU�?      �?        ��y��y�?�a�a�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?        �q�q�?��8��8�?      �?      �?�������?�?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        &���^B�?h/�����?      �?      �?]t�E�?F]t�E�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        r�q��?�q�q�?              �?�������?UUUUUU�?              �?      �?        ------�?�������?      �?      �?              �?      �?        �������?�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        к����?L�Ϻ��?�?xxxxxx�?�{a���?GX�i���?              �?      �?      �?              �?      �?      �?              �?      �?        ى�؉��?;�;��?(�����?�k(���?�������?�������?              �?      �?                      �?�������?ffffff�?t�E]t�?]t�E�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        9��8���?�q�q�?      �?              �?      �?              �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJUehG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       `                    �?|��;;��?�           8�@                                    @6kh�h��?�            �p@                                  �?PX�V|�?W            `a@                                 �;@      �?:             X@                                  �7@؇���X�?             5@                                  �6@�z�G��?             $@        ������������������������       �                     @               	                    �?      �?             @        ������������������������       �                      @        
                        ��m1@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@                                03�=@`2U0*��?.            �R@                                   �?�L���?            �B@                                03[:@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                  �B@Pa�	�?            �@@       ������������������������       �                     3@                                    �?@4և���?             ,@        ������������������������       �                     �?                                  �*@$�q-�?             *@                                  D@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     C@                                   @ qP��B�?            �E@        ������������������������       �                     �?        ������������������������       �                     E@                3                    �?�D}1o��?K             `@        !       2                 03�:@�T`�[k�?            �J@       "       #                   �+@��x_F-�?            �I@        ������������������������       �                      @        $       -                    �?>��C��?            �E@        %       *                    �?      �?             $@       &       '                 �%@���Q��?             @        ������������������������       �                      @        (       )                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        +       ,                   �-@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        .       /                 ���@6YE�t�?            �@@        ������������������������       �                     @        0       1                    �?��S�ۿ?             >@       ������������������������       �                     <@        ������������������������       �                      @        ������������������������       �                      @        4       Q                    �?,���y4�?/             S@       5       L                 ���1@�p ��?            �D@       6       C                   �7@     ��?             @@       7       B                    �?     ��?             0@       8       A                 �[$@���!pc�?	             &@       9       :                 ���@z�G�z�?             $@        ������������������������       �                     @        ;       @                 pF�!@�q�q�?             @       <       =                   �2@      �?             @        ������������������������       �                     �?        >       ?                   �6@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        D       E                   �&@      �?             0@       ������������������������       �                      @        F       G                    �?      �?              @        ������������������������       �                      @        H       I                 @3�/@�q�q�?             @        ������������������������       �                     �?        J       K                 �|�;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        M       P                 ���4@�����H�?             "@        N       O                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        R       ]                    @��R[s�?            �A@       S       V                    �?V�a�� �?             =@        T       U                 `f7@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        W       X                  `/@���}<S�?             7@        ������������������������       �                     �?        Y       \                    @���7�?             6@        Z       [                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             3@        ^       _                 ��T?@      �?             @        ������������������������       �                     @        ������������������������       �                     @        a       z                 �?�@2�Bo��?#           �{@        b       y                    �?X�Հ�+�?]            �`@       c       l                   �8@H*C�|F�?X             `@        d       g                    �?     ��?             @@        e       f                   �6@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        h       k                 ���@ 7���B�?             ;@        i       j                 ���@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     6@        m       n                  ��@`�E���?C            @X@        ������������������������       �        !            �G@        o       p                   �<@`2U0*��?"             I@        ������������������������       �                     .@        q       x                    �? >�֕�?            �A@        r       u                    �?�t����?             1@        s       t                 �|Y=@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        v       w                 X�I@ףp=
�?             $@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     @        {       �                   �;@N��c��?�            @s@        |       }                     �?䯦s#�?E            �Z@        ������������������������       �                     (@        ~       �                    �?p�v>��?=            �W@              �                    �?z�G�z�?"             I@        �       �                    (@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                     @:	��ʵ�?            �F@        �       �                    5@�IєX�?             1@       �       �                   �2@�C��2(�?             &@       ������������������������       �                     @        �       �                   �'@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    9@      �?             <@       �       �                 0S5 @���B���?             :@        �       �                   �3@X�Cc�?             ,@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     (@        ������������������������       �                      @        �       �                    �?8�A�0��?             F@        �       �                    �?z�G�z�?	             .@       �       �                    $@      �?             (@        ������������������������       �                     @        �       �                    7@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    #@l��[B��?             =@       �       �                   �C@�q�q�?             2@       �       �                    @$�q-�?	             *@       ������������������������       �                     $@        �       �                 ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?���!pc�?             &@        �       �                 ���)@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�#l��?�            @i@       �       �                     �?�,©T�?q            `f@        �       �                 ��9L@      �?-             Q@       �       �                   @J@r�����?#            �J@       �       �                   �G@����>�?            �B@       �       �                    �?     ��?             @@        �       �                 `f�A@      �?              @       �       �                 ��2>@      �?             @        ������������������������       �                      @        �       �                 X�lA@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �>@r�q��?             8@        �       �                 03:@���|���?             &@        ������������������������       �                     @        �       �                 �|�<@      �?              @        ������������������������       �                     �?        �       �                 03k:@և���X�?             @        ������������������������       �                     �?        �       �                 X��B@�q�q�?             @        �       �                 `fF<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �        	             *@        �       �                   �H@���Q��?             @        ������������������������       �                      @        �       �                   @I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             0@        �       �                 �|Y>@��S���?
             .@        ������������������������       �                     @        �       �                   �D@���|���?             &@        ������������������������       �                     @        �       �                    �?      �?              @       �       �                   @G@և���X�?             @        ������������������������       �                     @        �       �                   �H@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�@`�t�D7�?D            �[@        �       �                   �?@�eP*L��?             &@        ������������������������       �                      @        �       �                   �A@�q�q�?             "@        ������������������������       �z�G�z�?             @        ������������������������       �      �?             @        �       �                    �?�ڊ�e��??             Y@       �       �                    �?DE�SA_�?<            @X@       �       �                   �>@H0sE�d�?/            �R@        �       �                     @>A�F<�?             C@        �       �                   �'@�C��2(�?             &@        ������������������������       �                     @        �       �                 �|�=@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��) @�<ݚ�?             ;@        ������������������������       �                     ,@        �       �                 pf� @��
ц��?             *@        ������������������������       �                     @        �       �                 �|�=@�z�G��?             $@       �       �                   �<@�<ݚ�?             "@        ������������������������       �                     @        �       �                 ���"@�q�q�?             @        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @D@�?�|�?            �B@       ������������������������       �                     2@        �       �                   �'@�}�+r��?             3@        ������������������������       �                     &@        �       �                   �*@      �?              @        �       �                   �F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     6@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                 �ܭ2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                        �|Y>@�nkK�?             7@        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������|d�_Z�?�7s@K�?"=P9���?��1��?�&!��ȩ?��]tc�?      �?      �?�$I�$I�?۶m۶m�?333333�?ffffff�?              �?      �?      �?      �?              �?      �?              �?      �?                      �?{�G�z�?���Q��?L�Ϻ��?}���g�?      �?      �?              �?      �?        |���?|���?              �?�$I�$I�?n۶m۶�?              �?;�;��?�؉�؉�?�$I�$I�?۶m۶m�?      �?                      �?              �?              �?�}A_З?��}A�?      �?                      �?QW�uE�?W�uE]�?"5�x+��?���!5��?�?�������?              �?qG�w��?$�;��?      �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?      �?                      �?e�M6�d�?'�l��&�?      �?        �?�������?              �?      �?              �?        ������?����k�?dp>�c�?8��18�?      �?      �?      �?      �?t�E]t�?F]t�E�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?�������?333333�?      �?                      �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?        X|�W|��?PuPu�?��{a�?a���{�?UUUUUU�?UUUUUU�?              �?      �?        ӛ���7�?d!Y�B�?              �?�.�袋�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?V��K�?���݀��?t��:W�?Ũ�oS��?�7�yC�?�!oȫ?      �?      �?�������?�������?              �?      �?        	�%����?h/�����?�������?�������?      �?                      �?      �?        ?��W�?����?      �?        ���Q��?{�G�z�?      �?        ��+��+�?�A�A�?<<<<<<�?�?۶m۶m�?�$I�$I�?              �?      �?        �������?�������?۶m۶m�?�$I�$I�?      �?              �?              �?        �����?5�wL��?�����?�V�9�&�?              �?ڨ�l�w�?L� &W�?�������?�������?333333�?�������?              �?      �?        ��O��O�?l�l��?�?�?]t�E�?F]t�E�?      �?        �������?UUUUUU�?              �?      �?              �?              �?      �?��؉���?ى�؉��?%I�$I��?�m۶m��?              �?      �?              �?                      �?颋.���?/�袋.�?�������?�������?      �?      �?      �?        �������?333333�?              �?      �?              �?        GX�i���?���=��?UUUUUU�?UUUUUU�?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        F]t�E�?t�E]t�?      �?      �?              �?      �?              �?        �I��A��?��be�F�?~�Fu�?	��*�?      �?      �?Dj��V��?�V�9�&�?�u�)�Y�?���L�?      �?      �?      �?      �?      �?      �?              �?      �?      �?      �?                      �?      �?        �������?UUUUUU�?]t�E]�?F]t�E�?      �?              �?      �?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �?�������?      �?        F]t�E�?]t�E]�?              �?      �?      �?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?                      �?l��W���?Nq��$�?t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?��Q��?
ףp=
�?���_\�?����?��b�/��?O贁N�?������?Cy�5��?]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        9��8���?�q�q�?      �?        �;�;�?�؉�؉�?              �?ffffff�?333333�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?*�Y7�"�?к����?      �?        �5��P�?(�����?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�Mozӛ�?d!Y�B�?      �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�)�rhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       \                    �?"��p�?�           8�@                                   �?l��=���?�            p@                                   �?�:�^���?6            �V@                                  �?������?*             R@              
                 ��:3@P���Q�?             D@                                   �?"pc�
�?             &@       ������������������������       �                     @               	                 ���,@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     =@        ������������������������       �                     @@                                �|�:@�q�q�?             2@       ������������������������       �                     $@                                  @I@      �?              @                                    @؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               7                    �?hTe�E�?f            �d@              4                    L@z�09JX�?7            @X@              %                 `f$@t/*�?5            �W@               $                    ;@�\��N��?             3@              #                    �?�	j*D�?
             *@              "                 pf� @�q�q�?	             (@                               pf�@���!pc�?             &@        ������������������������       �                     @               !                   �9@      �?              @                                  �6@      �?             @                                   4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        &       3                    @HP�s��?&            �R@       '       2                    �?,N�_� �?%            �R@       (       1                    -@4��?�?             J@       )       *                 pF%@��hJ,�?             A@        ������������������������       �                     (@        +       0                    :@�GN�z�?	             6@        ,       /                 ��y)@r�q��?             @       -       .                 ��&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     0@        ������������������������       �                     2@        ������������������������       �                     6@        ������������������������       �                     �?        5       6                   �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        8       [                    @��(@��?/            �Q@       9       F                     @�2�,��?-            �P@        :       =                    6@�J�4�?             9@        ;       <                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        >       E                    �?���N8�?             5@       ?       @                   �E@�IєX�?             1@       ������������������������       �                     *@        A       D                   �F@      �?             @       B       C                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        G       N                   �1@����X�?             E@        H       I                     @և���X�?             ,@        ������������������������       �                      @        J       K                   -@      �?             (@        ������������������������       �                     @        L       M                 ��T?@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        O       Z                    �?؇���X�?             <@       P       Q                 �|Y=@��s����?             5@        ������������������������       �                     (@        R       W                     @X�<ݚ�?             "@       S       T                 �|Y>@      �?             @        ������������������������       �                      @        U       V                 03C3@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        X       Y                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ]       l                    *@ҔOl�?!           `|@        ^       c                    @`՟�G��?             ?@       _       b                    �?      �?             0@        `       a                 �y.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             *@        d       e                    �?�r����?	             .@        ������������������������       �                     @        f       k                    @r�q��?             (@       g       h                    �?���Q��?             @        ������������������������       �                      @        i       j                     @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        m       �                    �?v Og��?           pz@        n       �                     �?2lK����?2            @T@        o       z                  �}S@�G��l��?             E@       p       y                   �J@X�Cc�?             <@       q       x                 X�,@@ףp=
�?
             4@       r       w                    �?r�q��?             (@       s       t                 �|Y<@z�G�z�?             $@       ������������������������       �                     @        u       v                 �ܵ<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        {       �                    �?����X�?	             ,@       |                        p�w@���!pc�?             &@       }       ~                   �4@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 @�pX@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��K.@8�Z$���?            �C@       �       �                 ���@`Jj��?             ?@        ������������������������       �                     ,@        �       �                 ��� @�t����?             1@       �       �                    �?r�q��?	             (@       �       �                 �|Y=@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��d5@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�����H�?�            `u@       �       �                 ��$:@�a�^��?�            Pq@       �       �                     @\ ���?�            �m@        �       �                     �?�?�P�a�?(             N@        ������������������������       �                      @        �       �                   �*@���c���?"             J@       �       �                 �|�=@�T|n�q�?            �E@        �       �                    @      �?             8@        ������������������������       �                     @        �       �                 �|Y=@�z�G��?             4@       �       �                   �'@      �?             0@        �       �                    5@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �       �                   @D@�}�+r��?             3@       ������������������������       �        	             (@        �       �                   @G@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�n���k�?o             f@       �       �                 `�X#@p}"����?n            �e@       �       �                 ���"@`1�=7q�?d            �c@       �       �                   @@@�O��e�?^            �b@       �       �                 �Y�@�C��2(�?I            @^@        �       �                    �?h�����?             <@        ������������������������       �                      @        �       �                   �8@P���Q�?	             4@       �       �                 ���@�C��2(�?             &@        �       �                 ���@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?��r
'��?<            @W@        �       �                 �|Y=@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �>@������?5            �T@       �       �                 ��) @Х-��ٹ?1            �R@       �       �                 �?$@      �?*             P@        �       �                 �|�;@ףp=
�?             $@       ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                   �1@@3����?%             K@        ������������������������       �                     �?        ������������������������       �        $            �J@        �       �                 �|Y=@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        �       �                   �@և���X�?             @        ������������������������       �                      @        �       �                   �?@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     =@        �       �                 �|�=@����X�?             @       ������������������������       �                     @        �       �                   �?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             2@        ������������������������       �                      @        �       �                   �;@���Q��?             D@        ������������������������       �                      @        �       �                      @p�ݯ��?             C@       �       �                   �Q@h+�v:�?             A@       �       �                   �J@���|���?            �@@       �       �                    �?�f7�z�?             =@       �       �                   �G@և���X�?             <@       �       �                   �B@�q�q�?             8@       �       �                 03k:@�n_Y�K�?	             *@        ������������������������       �                     @        �       �                   @=@      �?             $@        �       �                 �|�?@      �?             @        ������������������������       �                      @        �       �                 `f�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 X�,C@�q�q�?             @       �       �                   @>@z�G�z�?             @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��9L@��ɉ�?*            @P@       ������������������������       �        #             M@        �       �                 `f�N@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @       �       �                 ��#[@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������J54v��?l�����?�`�`�`�?�'�'�'�?l�l��?}�'}�'�?�q�q�?�q�q�?�������?ffffff�?F]t�E�?/�袋.�?              �?�������?333333�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?۶m۶m�?�$I�$I�?              �?      �?                      �?�Ӛ��?@:�2	v�?W?���?:*����?W�+���?�;����?y�5���?�5��P�?;�;��?vb'vb'�?UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?              �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?                      �?      �?        {�G�z�?q=
ףp�?���L�?h�`�|��?ى�؉��?�N��N��?�������?KKKKKK�?              �?]t�E�?�袋.��?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?              �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?����?��+��+�?o�Wc"=�?"=P9���?{�G�z�?�z�G��?      �?      �?      �?                      �?�a�a�?��y��y�?�?�?              �?      �?      �?      �?      �?              �?      �?                      �?              �?�m۶m��?�$I�$I�?۶m۶m�?�$I�$I�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?z��y���?�a�a�?      �?        r�q��?�q�q�?      �?      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        z\��W&�?�$�f�?�s�9��?�1�c��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�?      �?        �������?UUUUUU�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ��X���?P$�Ҽ��?��a�2��?�<ݚ�?��y��y�?1�0��?�m۶m��?%I�$I��?�������?�������?UUUUUU�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        �m۶m��?�$I�$I�?F]t�E�?t�E]t�?�q�q�?�q�q�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?;�;��?���{��?�B!��?      �?        <<<<<<�?�?�������?UUUUUU�?/�袋.�?F]t�E�?              �?      �?              �?              �?              �?      �?              �?      �?        �q�q�?�q�q�?��U��?�'�3���?�O�%�L�?����v��?DDDDDD�?�����ݽ?      �?        ;�;��?�;�;�?���)k��?6eMYS��?      �?      �?      �?        ffffff�?333333�?      �?      �?�m۶m��?�$I�$I�?              �?      �?              �?                      �?�5��P�?(�����?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?        a��S��?��i�`Ͳ?ĦҐs��?��jyc�?b��x�Y�?�\�:�2�?�t�@��?ƒ_,�Ų?]t�E�?F]t�E�?�m۶m��?�$I�$I�?      �?        ffffff�?�������?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?              �?        �<��#��?�n�ᆻ?/�袋.�?F]t�E�?              �?      �?        �|����?������?K~��K�?O贁N�?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?���Kh�?h/�����?              �?      �?        /�袋.�?F]t�E�?      �?                      �?۶m۶m�?�$I�$I�?              �?333333�?�������?              �?      �?              �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        333333�?�������?              �?^Cy�5�?Cy�5��?�������?xxxxxx�?]t�E]�?F]t�E�?O#,�4��?a���{�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?ى�؉��?;�;��?              �?      �?      �?      �?      �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?              �?      �?              �?                      �?      �?              �?                      �?      �?      �?      �?                      �??�?��? �����?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJX"4qhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMAhjh))��}�(h,h/h0MA��h2h3h4hph<�h=Kub������       f                 ���"@|��;;��?�           8�@               !                    �?J��ԛ�?�            �m@                                    �?�萻/#�?-            �P@                                  �?8�A�0��?,            �P@        ������������������������       �                     3@                                ���@t/*�?            �G@                                03S@��S�ۿ?             .@        ������������������������       �                      @        	       
                 �|�9@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@                                   �?     ��?             @@                                  @8@������?             .@        ������������������������       �                      @                                �|�=@8�Z$���?
             *@                                 �<@      �?              @        ������������������������       �                      @                                  @@�q�q�?             @       ������������������������       ��q�q�?             @                                �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                ���@@�0�!��?             1@        ������������������������       �                     @                                �|Y=@���!pc�?             &@        ������������������������       �                     �?                                X�I@z�G�z�?             $@                               ��(@�<ݚ�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        "       e                    �?x�ۈp�?o            `e@       #       d                   @D@<���i�?n            @e@       $       5                    �?      �?d             c@        %       .                 P�@��
ц��?             *@       &       -                    �?����X�?             @       '       ,                 �|�;@���Q��?             @       (       )                 pf�@      �?             @        ������������������������       �                      @        *       +                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        /       4                 `�X!@�q�q�?             @       0       3                    �?z�G�z�?             @       1       2                   �8@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        6       7                     @��˥W1�?Y            `a@        ������������������������       �        	             *@        8       c                    �?�����?P            �_@       9       b                    �?������?O            �^@       :       _                    �?�D�d@6�?M            �]@       ;       L                 �?�@t��%�?I            �\@       <       =                   �7@0�,���?,            �P@        ������������������������       �                     3@        >       K                 �?$@ �q�q�?              H@       ?       F                 ���@ 	��p�?             =@       @       E                   �8@�nkK�?             7@        A       D                 `fF@      �?             @       B       C                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        G       H                 �|�;@r�q��?             @        ������������������������       �                      @        I       J                 �|Y>@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     3@        M       P                 @3�@     ��?             H@        N       O                   �A@�n_Y�K�?             *@       ������������������������       �                     @        ������������������������       �����X�?             @        Q       X                 ��i @(N:!���?            �A@       R       U                   �3@؇���X�?             5@        S       T                   �1@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �      �?              @        V       W                 ��) @      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?        Y       Z                 pf� @@4և���?             ,@        ������������������������       �                     @        [       \                    8@�C��2(�?             &@        ������������������������       �                     @        ]       ^                    <@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        `       a                 P�@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             2@        ������������������������       �                     �?        g       *                @�:R@��;�4��?#           �}@       h       #                   @(옄��?�            �y@       i       �                     @�7 ����?�            �w@       j       �                    �?�Nj���?�            �o@        k       r                     �?�����H�?<             [@        l       q                    �? �q�q�?             8@        m       p                    �?؇���X�?             @        n       o                   �B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        s       �                    �?H��?"�?0             U@        t       {                   @B@�㙢�c�?             G@       u       z                   �9@(;L]n�?             >@        v       y                    �?$�q-�?             *@        w       x                   �6@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             1@        |       �                   �*@     ��?             0@       }       �                   �'@��
ц��?             *@        ~                          �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    D@      �?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�˹�m��?             C@        ������������������������       �                     @        �       �                    6@     ��?             @@        �       �                   �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��S�ۿ?             >@       �       �                   �E@�>����?             ;@       ������������������������       �                     3@        �       �                   �8@      �?              @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�c�Α�?Y             b@       �       �                     �?��ٌ���?X            �a@        �       �                    �?�J�T�?'            �Q@       �       �                    �?`�(c�?            �H@        �       �                 p�i@@�E��ӭ�?             2@       �       �                 ���=@�eP*L��?             &@        ������������������������       �                     @        �       �                  Y>@      �?              @        ������������������������       �                     @        �       �                 X�lA@���Q��?             @        ������������������������       �                      @        �       �                  �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �;@`՟�G��?             ?@        ������������������������       �                      @        �       �                    R@�f7�z�?             =@       �       �                   �>@��}*_��?             ;@       �       �                    M@      �?
             0@       �       �                 ��<:@�θ�?             *@        ������������������������       �                     �?        �       �                 `f�;@r�q��?             (@        ������������������������       �                     @        �       �                 X��B@����X�?             @        ������������������������       �                     @        �       �                   �=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                      @        �       �                 �5L@"pc�
�?	             6@       �       �                 `�iJ@      �?             0@        �       �                  x#J@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 0��M@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    #@�q�q�?1             R@        ������������������������       �                     $@        �       �                    �?6uH���?,             O@       �       �                    �?�����H�?            �F@       �       �                    �?�Ra����?             F@        ������������������������       �                     �?        �       �                    @@X�EQ]N�?            �E@       �       �                    &@���7�?             6@        �       �                    5@      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        
             ,@        �       �                   @A@��s����?             5@        ������������������������       �                     @        �       �                    F@�X�<ݺ?             2@        �       �                   �3@      �?              @        �       �                   @D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                      @        �                          @v�2t5�?N            �^@       �       �                    �?f=UBS�?I            @]@        �       �                    �?`�(c�?             �H@        �       �                    �?���!pc�?             6@       �       �                 �|Y=@      �?	             0@       �       �                    �?"pc�
�?             &@        ������������������������       �                     @        �       �                    '@�q�q�?             @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                  S�2@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?|��?���?             ;@        �       �                    �?      �?              @       �       �                    4@z�G�z�?             @        ������������������������       �                     @        �       �                   P&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �@@p�ݯ��?             3@       �       �                    �?������?             .@       �       �                    �?�	j*D�?
             *@        �       �                 03�0@�q�q�?             @       �       �                 ���)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    0@����X�?             @        ������������������������       �                     �?        �       �                 `fv1@r�q��?             @        ������������������������       �                     @        �       �                 `fV6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 `f�/@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                               �T)D@�t����?)             Q@                                �?�w��@�?&            �O@                                 �?�<ݚ�?             "@                                3@���Q��?             @        ������������������������       �                      @                                 �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        	      
                   )@r�q��?!             K@        ������������������������       �                     @                              �|�=@Hm_!'1�?            �H@                                �?      �?             @@        ������������������������       �                      @                              `�X#@ �q�q�?             8@                                �<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@                              ���'@@�0�!��?	             1@                                �?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@                              �|�;@z�G�z�?             @        ������������������������       �                     @                              �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 @r�q��?             @        ������������������������       �                     @              "                   @�q�q�?             @              !                ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        $      %                ��T?@�}�+r��?             C@       ������������������������       �                     8@        &      )                   @؇���X�?	             ,@        '      (                   �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        +      ,                   �?0B��D�?)            �M@       ������������������������       �                    �B@        -      .                 �}S@�X����?             6@        ������������������������       �                      @        /      8                   �?      �?             4@       0      1                Ј�V@z�G�z�?             $@        ������������������������       �                     @        2      3                   �?���Q��?             @        ������������������������       �                      @        4      7                   �?�q�q�?             @       5      6                  �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        9      :                0�X@�z�G��?             $@        ������������������������       �                     �?        ;      <                   6@�<ݚ�?             "@        ������������������������       �                     �?        =      @                   �?      �?              @       >      ?                   �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MAKK��h2h3h4hVh<�h=Kub������������|d�_Z�?�7s@K�?�ԋ�ԋ�?�����?ï�Dz��?z�rv��?颋.���?/�袋.�?              �?�;����?W�+���?�������?�?      �?        �؉�؉�?;�;��?              �?      �?              �?      �?wwwwww�?�?              �?;�;��?;�;��?      �?      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        ZZZZZZ�?�������?      �?        F]t�E�?t�E]t�?              �?�������?�������?9��8���?�q�q�?      �?      �?      �?              �?                      �?�w�A�?�A|�?llllll�?�������?      �?      �?�؉�؉�?�;�;�?�$I�$I�?�m۶m��?�������?333333�?      �?      �?              �?      �?      �?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?ۻ��<�?'!����?      �?        =��<���?�a�a�?�|����?������?}��|���?���й?�(�j��?�q�.�|�?Ez�rv�?g��1��?      �?        �������?UUUUUU�?������?�{a���?�Mozӛ�?d!Y�B�?      �?      �?      �?      �?      �?                      �?      �?              �?        �������?UUUUUU�?      �?              �?      �?      �?      �?      �?              �?              �?      �?;�;��?ى�؉��?      �?        �$I�$I�?�m۶m��?|�W|�W�?�A�A�?۶m۶m�?�$I�$I�?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?      �?        ]t�E�?F]t�E�?      �?        �������?�������?              �?      �?              �?      �?      �?                      �?      �?              �?              �?                      �?l��	�<�?(��Æ�?���,d�?ӛ���7�?�+���?�٨�l��?X_ʘ�?�SqК3�?�q�q�?�q�q�?UUUUUU�?�������?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?1�0��?�<��<��?d!Y�B�?�7��Mo�?�?�������?;�;��?�؉�؉�?�������?�������?              �?      �?                      �?              �?      �?      �?�;�;�?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?              �?^Cy�5�?��P^Cy�?              �?      �?      �?      �?      �?              �?      �?        �?�������?h/�����?�Kh/��?              �?      �?      �?              �?      �?      �?      �?                      �?              �?5�rO#,�?�{a���?	�g��?�U0K��?H���@��?p�z2~��?������?4և����?�q�q�?r�q��?t�E]t�?]t�E�?      �?              �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �1�c��?�s�9��?              �?O#,�4��?a���{�?_B{	�%�?B{	�%��?      �?      �?�؉�؉�?ى�؉��?      �?        UUUUUU�?�������?              �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?/�袋.�?F]t�E�?      �?      �?�������?�������?      �?                      �?      �?              �?      �?              �?      �?        UUUUUU�?�������?              �?k���Zk�?��RJ)��?�q�q�?�q�q�?]t�E]�?]t�E�?      �?        w�qG�?qG�wĽ?�.�袋�?F]t�E�?      �?      �?      �?      �?      �?              �?        z��y���?�a�a�?              �?��8��8�?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?              �?                      �?��+Q��?�ڕ�]��?2%S2%S�?��Y��Y�?4և����?������?t�E]t�?F]t�E�?      �?      �?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?                      �?              �?	�%����?{	�%���?      �?      �?�������?�������?              �?      �?      �?      �?                      �?              �?^Cy�5�?Cy�5��?wwwwww�?�?vb'vb'�?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?�������?�������?�}��}��?AA�?�q�q�?9��8���?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?UUUUUU�?              �?Y�Cc�?9/���?      �?      �?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        ZZZZZZ�?�������?      �?      �?              �?      �?              �?        �������?�������?              �?      �?      �?      �?                      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �5��P�?(�����?      �?        ۶m۶m�?�$I�$I�?333333�?�������?      �?                      �?      �?        ��}ylE�?�A�I��?              �?�E]t��?]t�E]�?              �?      �?      �?�������?�������?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?ffffff�?333333�?              �?9��8���?�q�q�?              �?      �?      �?�������?UUUUUU�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ;�3whG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       n                     @�����?�           8�@                                   �?bf@����?�            �s@                                   �? �#�Ѵ�?Y             `@                                  �?@4և���?:             U@                                   �?�}�+r��?             C@                               03�=@$�q-�?             :@               
                    �?      �?             @              	                     �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                     (@                                   L@���}<S�?#             G@                                 �;@��S�ۿ?"            �F@                                    �?z�G�z�?             $@        ������������������������       �                     �?                                  �7@�<ݚ�?             "@                                 �6@���Q��?             @        ������������������������       �                      @                                  �'@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                  �E@��?^�k�?            �A@       ������������������������       �                     =@                                   �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �F@                '                   �1@����c��?n            `g@        !       &                    �?$�q-�?             *@        "       #                     �?      �?             @        ������������������������       �                      @        $       %                 ���?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        (       A                 ��D:@�s��9n�?h            �e@        )       @                    �?�:�^���?0            �S@       *       ?                    F@ ����?)            @P@       +       >                   �D@^�!~X�?!            �J@       ,       =                   @A@ i���t�?            �H@       -       <                    @@�ݜ�?            �C@       .       1                    5@�L���?            �B@        /       0                    &@z�G�z�?             $@        ������������������������       ����Q��?             @        ������������������������       �                     @        2       3                     �? 7���B�?             ;@        ������������������������       �                     @        4       5                 �|Y=@ �q�q�?             8@       ������������������������       �        
             0@        6       7                    @      �?              @        ������������������������       �                     @        8       9                    �?z�G�z�?             @        ������������������������       �                     �?        :       ;                 �|�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �      �?             @        ������������������������       �                     (@        ������������������������       �                     *@        B       m                   �J@     ��?8             X@       C       l                     �?�Jhu4��?+            @R@       D       k                    �?     ��?$             P@       E       R                  �>@�g�y��?#             O@        F       Q                    @@��+7��?             7@       G       H                    <@��
ц��?             *@        ������������������������       �                     @        I       P                   @>@�q�q�?             "@       J       K                    �?؇���X�?             @        ������������������������       �                      @        L       M                 `fF<@z�G�z�?             @        ������������������������       �                      @        N       O                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        S       X                 �|Y<@�q�q�?            �C@        T       W                    �?؇���X�?             @       U       V                 �U�X@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        Y       Z                 �|Y>@     ��?             @@        ������������������������       �                     &@        [       j                   �H@�q�q�?             5@       \       i                   �G@j���� �?             1@       ]       h                    �?����X�?             ,@       ^       g                    �?���Q��?             $@       _       f                   �E@X�<ݚ�?             "@       `       a                   �A@և���X�?             @        ������������������������       �                      @        b       c                    �?���Q��?             @        ������������������������       �                      @        d       e                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     7@        o       �                 P��%@�o6�
�?�            �x@       p       q                 ���@"pc�
�?�            �o@        ������������������������       �                     7@        r       �                    �?z�G�z�?�            �l@        s       |                 �|Y=@�99lMt�?            �C@       t       {                    �?�\��N��?             3@       u       z                 03�!@�θ�?
             *@       v       w                 �?@�C��2(�?	             &@       ������������������������       �                     @        x       y                   �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        }       ~                    �?      �?
             4@       ������������������������       �                     (@               �                 �|Y>@      �?              @        ������������������������       �                     @        �       �                    C@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��@p^�AL�?x            �g@        ������������������������       �                     �?        �       �                ��k @�KM�]�?w            �g@        ������������������������       �                      @        �       �                   @@@��8��)�?v            �g@       �       �                 ���"@�	L �F�?b            `c@       �       �                  ��@ܷ��?��?[             b@        �       �                 �Y�@ 7���B�?             ;@        �       �                    �?@4և���?
             ,@       �       �                 ���@$�q-�?	             *@       ������������������������       �                     @        �       �                   @8@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             *@        �       �                    �?�^����?G            �]@        ������������������������       �                     @        �       �                    �?���5��?E            �\@        �       �                 ��(@z�G�z�?
             .@       �       �                    �?d}h���?	             ,@       �       �                 �|Y=@���!pc�?             &@        ������������������������       �                     �?        ������������������������       �z�G�z�?             $@        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�����H�?;            �X@       �       �                 �|�>@�W�{�5�?9            �W@       �       �                 �?$@|)����?7            �V@        �       �                 �|�;@      �?             (@       ������������������������       �                     @        ������������������������       ����Q��?             @        �       �                 �?�@86��Z�?1            �S@        ������������������������       �                    �D@        �       �                   �4@�?�'�@�?             C@        �       �                 0S5 @���!pc�?	             &@        �       �                   �2@���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �9@�>����?             ;@        ������������������������       �                     $@        �       �                    <@�t����?             1@        ������������������������       �                     �?        �       �                 ��) @      �?
             0@       ������������������������       �                     (@        �       �                 pf� @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 P�@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���#@�z�G��?             $@       �       �                   �<@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �@@        �       �                    �?���W�?]            �a@        �       �                 ��Y7@ꮃG��?.            @Q@       �       �                    @Z�K�D��?            �G@        �       �                 ��*4@��S�ۿ?	             .@       ������������������������       �                     &@        �       �                 �̌5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @      �?             @@       �       �                    5@�g�y��?             ?@        �       �                    �?      �?             (@       �       �                    �?      �?              @        �       �                   �-@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��.@p�ݯ��?             3@        �       �                 �|Y<@����X�?             @        ������������������������       �                     �?        �       �                 ��*@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?	             (@        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                     @      �?             @       �       �                 ��1@�q�q�?             @       �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?"pc�
�?             6@        ������������������������       �                     �?        �       �                    @؇���X�?             5@        ������������������������       �                      @        �       �                    �?�}�+r��?             3@        ������������������������       �                     �?        �       �                 X��@@�X�<ݺ?             2@       ������������������������       �        
             .@        �       �                    @�q�q�?             @        ������������������������       �                     �?        �       �                 pf�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    *@z�z�7��?/            @R@        �       �                    @��H�}�?             9@        �       �                    �?�����H�?             "@       ������������������������       �                     @        �       �                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `f68@      �?             0@        ������������������������       �                     @        �       �                 ��A>@z�G�z�?             $@       ������������������������       �                     @        �       �                 pf�C@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �                          �?�8��8��?             H@                                  �?؇���X�?             @                             �|Y<@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?��p\�?            �D@                              �T)D@     ��?
             0@       ������������������������       �                     &@              	                   ;@���Q��?             @        ������������������������       �                      @        
                      �|�>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     9@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�����������������?��܍��?T:�g *�?��&��j�?�}A_Ч?�/����?�$I�$I�?n۶m۶�?(�����?�5��P�?;�;��?�؉�؉�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?d!Y�B�?ӛ���7�?�?�������?�������?�������?              �?�q�q�?9��8���?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�A�A�?_�_��?              �?UUUUUU�?�������?              �?      �?              �?                      �?�W@�n��?�P9"��?;�;��?�؉�؉�?      �?      �?              �?      �?      �?      �?                      �?              �?^ ��2�?�~�u�7�?� � �?�o��o��?�ȍ�ȍ�?�����?�}�	��?�	�[���?/�����?����X�?\��[���?�i�i�?}���g�?L�Ϻ��?�������?�������?333333�?�������?      �?        	�%����?h/�����?      �?        �������?UUUUUU�?      �?              �?      �?      �?        �������?�������?      �?              �?      �?              �?      �?                      �?      �?              �?      �?      �?              �?              �?      �?�-[�l��?ҤI�&M�?      �?      �?�B!��?��{���?Y�B��?zӛ����?�؉�؉�?�;�;�?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?�������?ZZZZZZ�?�m۶m��?�$I�$I�?333333�?�������?r�q��?�q�q�?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?                      �?      �?              �?              �?              �?        �}z)@w�?	Z�"�?/�袋.�?F]t�E�?      �?        �������?�������?�o��o��?5H�4H��?�5��P�?y�5���?�؉�؉�?ى�؉��?F]t�E�?]t�E�?              �?�������?�������?      �?                      �?      �?              �?              �?      �?              �?      �?      �?      �?              �?      �?              �?      �?        i�O{�?��)_�%�?              �?�k(���?(�����?              �?�Q�٨��?br1���?I��īH�?��ۡ��?��=���?a���{�?	�%����?h/�����?n۶m۶�?�$I�$I�?�؉�؉�?;�;��?      �?        �������?UUUUUU�?              �?      �?              �?              �?        u_[4�?W'u_�?      �?        �}��?��Gp�?�������?�������?I�$I�$�?۶m۶m�?F]t�E�?t�E]t�?              �?�������?�������?      �?              �?        �q�q�?�q�q�?�ĩ�sK�?Fڱa��?��/��/�?h�h��?      �?      �?      �?        �������?333333�?�Z܄��?h *�3�?      �?        ������?y�5���?F]t�E�?t�E]t�?�������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        �Kh/��?h/�����?      �?        <<<<<<�?�?              �?      �?      �?      �?              �?      �?              �?      �?              �?      �?              �?      �?              �?        ffffff�?333333�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ��9�h�?ܥ���.�?s��\;�?�%~F��?]AL� &�?R�٨�l�?�?�������?              �?      �?      �?      �?                      �?      �?      �?�B!��?��{���?      �?      �?      �?      �?�������?333333�?      �?                      �?      �?              �?        Cy�5��?^Cy�5�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?�$I�$I�?�m۶m��?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?              �?              �?/�袋.�?F]t�E�?              �?۶m۶m�?�$I�$I�?              �?�5��P�?(�����?      �?        ��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ҤI�&M�?�lٲe��?{�G�z�?
ףp=
�?�q�q�?�q�q�?      �?              �?      �?              �?      �?              �?      �?              �?�������?�������?      �?        333333�?�������?              �?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?                      �?      �?        �]�ڕ��?��+Q��?      �?      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�3hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM)hjh))��}�(h,h/h0M)��h2h3h4hph<�h=Kub������       �                     @�E	�rQ�?�           8�@                                  �1@)b���?�            t@                                   �?HP�s��?             9@       ������������������������       �        	             4@                                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @               {                    �?�hP���?�            �r@       	       J                     �?�AS���?�            `n@       
                           �?X�<ݚ�?T            �`@                                  �H@4��?�?              J@       ������������������������       �                     D@                                   �?�q�q�?             (@                                  �?X�<ݚ�?             "@                                  K@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               I                 ��v@j����?4            �T@              "                    �?     ��?3             T@                                  �8@��
ц��?             :@        ������������������������       �                     @               !                   �H@p�ݯ��?             3@                               �|Y<@؇���X�?
             ,@        ������������������������       �                     @                                  �>@����X�?             @                                �ܵ<@�q�q�?             @        ������������������������       �                     �?                                ��2>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        #       <                   �G@����|e�?#             K@       $       5                    �?r�q��?             E@       %       (                 �|�<@�<ݚ�?             ;@        &       '                 `f�D@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        )       .                   �@@r�q��?             8@       *       -                   �>@�IєX�?	             1@        +       ,                   �1@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        /       0                   �9@և���X�?             @        ������������������������       �                      @        1       2                    D@���Q��?             @        ������������������������       �                      @        3       4                  I>@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        6       7                   �C@��S�ۿ?             .@        ������������������������       �                     @        8       ;                 0�nL@      �?              @        9       :                  x#J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        =       @                 `fF<@      �?             (@        >       ?                    J@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        A       D                   �I@����X�?             @        B       C                 ���W@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        E       F                   �J@z�G�z�?             @        ������������������������       �                     @        G       H                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        K       d                    �?�Sb(�	�?G             [@        L       c                    L@�MI8d�?            �B@       M       T                   �;@4?,R��?             B@        N       S                   �7@���!pc�?             &@       O       P                    �?      �?             @        ������������������������       �                      @        Q       R                 ��m1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        U       `                    9@HP�s��?             9@       V       W                 ��Y)@�}�+r��?             3@        ������������������������       �                     @        X       _                    �?$�q-�?
             *@       Y       Z                   �B@�8��8��?	             (@       ������������������������       �                     @        [       ^                   �,@z�G�z�?             @        \       ]                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        a       b                    D@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        e       t                   @D@����Q8�?+            �Q@       f       s                 ��,@h㱪��?!            �K@       g       l                    4@���N8�?             E@        h       i                   �2@      �?              @       ������������������������       �                     @        j       k                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        m       n                 �|Y=@г�wY;�?             A@        ������������������������       �        
             .@        o       p                   �'@�}�+r��?             3@       ������������������������       �                     (@        q       r                 �|�=@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        u       z                   �*@      �?
             0@       v       w                 `f�)@�<ݚ�?             "@        ������������������������       �                     @        x       y                    G@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        |       �                   �L@r�z-��?             �J@       }       �                    �?�<ݚ�?            �F@       ~       �                  D�Y@R�}e�.�?             :@              �                    �?     ��?             0@        �       �                    �?և���X�?             @        ������������������������       �                     @        �       �                 `��Q@      �?             @       �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�S����?             3@       ������������������������       �        	             0@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?f]��U�?�            `x@       �       �                    �?�%�\�@�?�            �q@        �       �                    �?�#}7��?)            �P@        �       �                    �?4?,R��?             B@       �       �                    �?�8��8��?             8@        ������������������������       �                     �?        �       �                 ���@���}<S�?             7@        ������������������������       �                      @        ������������������������       �                     5@        �       �                    �?      �?             (@        �       �                 �|Y6@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   @D@�P�*�?             ?@       �       �                 �|Y>@П[;U��?             =@       �       �                    �?�n_Y�K�?             :@       �       �                  sW@���Q��?             4@        �       �                 pf�@      �?              @       ������������������������       �                     @        �       �                    4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��&@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                 ���)@�q�q�?             @       ������������������������       �                     @        �       �                 03�0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                  ��@�~i��?�            @k@        �       �                   @4@ �Jj�G�?(            �K@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        $            �I@        �       �                 �T)D@�Ǐ�?f            `d@       �       �                    �?�v,D�?c            �c@        �       �                 �|Y=@$�q-�?             *@        �       �                   �;@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?\-��p�?\             b@       �       �                    �?8�Z$���?R            @`@        �       �                 ��(@z�G�z�?
             .@       �       �                 �|Y=@d}h���?	             ,@        ������������������������       �                     �?        �       �                 X��A@8�Z$���?             *@       ������������������������       �"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���#@V�n���?H            �\@       �       �                 �?�@�v�G���?@            �Y@        �       �                 �|�<@��-�=��?            �C@       ������������������������       �                     7@        �       �                   @@@      �?
             0@       �       �                    ?@�	j*D�?             *@       �       �                  sW@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                   �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@     ��?'             P@        �       �                   �A@      �?              @       �       �                    :@����X�?             @        ������������������������       �                      @        �       �                   �?@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        �       �                   �0@�>4և��?              L@        �       �                 �̌!@�q�q�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        �       �                 ���"@H%u��?             I@       �       �                   �3@��(\���?             D@        �       �                    2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        �       �                   �:@ >�֕�?            �A@        ������������������������       �                     0@        �       �                 �|Y<@�KM�]�?             3@        ������������������������       �                     �?        �       �                 ��) @�X�<ݺ?             2@       ������������������������       �        	             ,@        �       �                 ��y @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�=@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �        
             .@        �       �                    ;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �                          �?n�����?<            @Z@        �       �                    @8����?             7@        ������������������������       �                     @        �       �                    �?     ��?
             0@       �       �                   �7@�q�q�?             "@        ������������������������       �                     @        �       �                    �?      �?             @       �       �                 �|Y=@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                 �2@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @              (                   @���� �?.            �T@                                �?�(�Tw��?+            �S@        ������������������������       �                     "@                                 �?4�	~���?'            @Q@                                �?����>�?            �B@                                �;@�q�q�?	             (@       	      
                @3�2@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                 @z�G�z�?             9@                                @���N8�?
             5@                              �̼6@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@                              ��T?@�q�q�?             "@                                ,@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @              '                   @      �?             @@                                @�f7�z�?             =@                                 @�C��2(�?             &@        ������������������������       �                     @                                 @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @              &                   @�����H�?             2@              %                   �?"pc�
�?             &@       !      "                P��)@�<ݚ�?             "@        ������������������������       �                     �?        #      $                   )@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M)KK��h2h3h4hVh<�h=Kub�������������JP���?7j_Q��?��4>2��?����f��?{�G�z�?q=
ףp�?              �?�������?333333�?      �?                      �?0E>�S�?�u�)�Y�?W�$﯃�?QA�!���?�q�q�?r�q��?ى�؉��?�N��N��?              �?�������?�������?r�q��?�q�q�?�������?UUUUUU�?      �?                      �?              �?              �?f�@	o4�?4u~�!��?      �?      �?�;�;�?�؉�؉�?      �?        Cy�5��?^Cy�5�?�$I�$I�?۶m۶m�?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        ����K�?	�%����?�������?UUUUUU�?9��8���?�q�q�?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?�?�?�������?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        �������?�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?�������?�������?              �?      �?        �$I�$I�?�m۶m��?      �?      �?      �?                      �?�������?�������?              �?      �?      �?      �?                      �?              �?�Kh/��?�Kh/���?L�Ϻ��?��L���?r�q��?�8��8��?t�E]t�?F]t�E�?      �?      �?              �?      �?      �?              �?      �?                      �?{�G�z�?q=
ףp�?(�����?�5��P�?              �?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?UUUUUU�?�������?              �?      �?              �?        O�o�z2�?��Vج?־a���?��)A��?��y��y�?�a�a�?      �?      �?      �?              �?      �?              �?      �?        �?�?      �?        �5��P�?(�����?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?              �?      �?9��8���?�q�q�?      �?        333333�?�������?              �?      �?              �?        �琚`��?����!�?�q�q�?9��8���?�;�;�?'vb'vb�?      �?      �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?              �?      �?              �?                      �?�������?333333�?              �?      �?        ^Cy�5�?(������?              �?      �?              �?        �tM�tM�?QeQe�?ׅ'�j]�?��aoT��?���[��?~5&��?r�q��?�8��8��?UUUUUU�?UUUUUU�?              �?d!Y�B�?ӛ���7�?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?�RJ)���?�Zk����?�{a���?��=���?;�;��?ى�؉��?333333�?�������?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ��w� z�?��A��.�?k߰�k�?��)A��?      �?      �?              �?      �?              �?        ]w��|�?�"���?~W��0��?�ґ=�?�؉�؉�?;�;��?      �?      �?      �?                      �?      �?        a����?�{a���?;�;��?;�;��?�������?�������?I�$I�$�?۶m۶m�?              �?;�;��?;�;��?/�袋.�?F]t�E�?      �?              �?        ���9E�?/�|���?C���?��O �?}˷|˷�?�A�A�?      �?              �?      �?vb'vb'�?;�;��?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?             ��?      �?      �?      �?�m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?      �?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?�������?�������?      �?        )\���(�?���Q��?�������?333333�?�������?�������?      �?              �?      �?��+��+�?�A�A�?      �?        �k(���?(�����?              �?��8��8�?�q�q�?      �?              �?      �?              �?      �?        ffffff�?333333�?      �?                      �?      �?              �?        333333�?�������?              �?      �?        �Fk�Fk�?�r)�r)�?8��Moz�?d!Y�B�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?333333�?�������?              �?      �?                      �?�$I�$I�?۶m۶m�?      �?                      �?jW�v%j�?,Q��+�?�o��o��?� � �?      �?        ];0���?F��Q�g�?�u�)�Y�?���L�?�������?�������?UUUUUU�?�������?              �?      �?              �?        �������?�������?�a�a�?��y��y�?�������?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?              �?      �?              �?      �?O#,�4��?a���{�?F]t�E�?]t�E�?              �?�������?�������?      �?                      �?�q�q�?�q�q�?/�袋.�?F]t�E�?9��8���?�q�q�?              �?      �?      �?              �?      �?              �?              �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ� �NhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       T                    �?�t����?�           8�@               Q                 p�H@�桐-�?�            @p@                                  �?�%�aW	�?t            �f@                                   �?���*�?%             N@                                  �?Du9iH��?            �E@       ������������������������       �                     :@                                   �?@�0�!��?             1@              	                     @�q�q�?             "@        ������������������������       �                     @        
                        �|Y6@      �?             @                                 �-@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                   �?��.k���?             1@                                  �?���Q��?	             .@                               `�@1@�eP*L��?             &@                                  �?      �?              @        ������������������������       �                     @                                �|Y=@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @               :                    �?�q�q�?O            �^@              1                    �?��X���?+            @Q@              .                 �|�=@�+e�X�?             I@              #                     @f���M�?             ?@               "                   �9@�C��2(�?             &@                !                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        $       +                   �@      �?             4@        %       *                 pff@z�G�z�?             $@        &       '                 ���@�q�q�?             @        ������������������������       �                     @        (       )                 �|Y:@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ,       -                    3@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        /       0                 ��n @�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        2       3                     @�}�+r��?             3@       ������������������������       �                     *@        4       5                    �?r�q��?             @        ������������������������       �                      @        6       7                    @      �?             @        ������������������������       �                      @        8       9                 ��l4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ;       L                    @|��?���?$             K@       <       C                     @X�<ݚ�?            �F@       =       B                    :@ �q�q�?             8@       >       ?                   �E@�X�<ݺ?             2@       ������������������������       �        
             0@        @       A                   �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        D       E                    #@�����?             5@        ������������������������       �                     �?        F       G                 ���.@P���Q�?             4@        ������������������������       �                     $@        H       K                 03�0@ףp=
�?             $@        I       J                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        M       N                    �?�����H�?             "@        ������������������������       �                     @        O       P                   �0@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        R       S                      @�g<a�?/            @S@       ������������������������       �        -            �R@        ������������������������       �                      @        U       �                  x#J@���{.��?,           0|@       V       q                 �?�@|D�]�|�?           �x@        W       p                    �?�?�0�!�?_             a@       X       ]                   @4@     8�?Y             `@        Y       Z                 �Y�@8�Z$���?             *@        ������������������������       �                     @        [       \                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ^       _                   �<@��x$�?Q            �\@        ������������������������       �                     <@        `       a                     @XB���?:            �U@        ������������������������       �                     $@        b       c                 ���@`<)�+�?4            @S@        ������������������������       �                    �@@        d       g                 �|Y=@t��ճC�?             F@        e       f                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        h       i                    �?������?            �D@        ������������������������       �                     @        j       o                   @@@ >�֕�?            �A@       k       n                   �@�>����?             ;@        l       m                    �?؇���X�?	             ,@       ������������������������       �$�q-�?             *@        ������������������������       �                     �?        ������������������������       �        
             *@        ������������������������       �                      @        ������������������������       �                      @        r       }                    @��3��?�            `p@        s       t                     @      �?	             (@        ������������������������       �                     @        u       x                    �?և���X�?             @        v       w                 03�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        y       |                     @      �?             @       z       {                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ~       �                    $@�L����?�            @o@               �                    @���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                 @3�@�d���?�             n@        �       �                   �9@�q�q�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �?@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        �       �                    �?��|��?�            @m@       �       �                    �?���?�             l@       �       �                 `fF:@���ZӼ�?�             i@       �       �                   �*@@݈g>h�?b             c@       �       �                    �?��8����?@             X@       �       �                   �3@Df/��?>            �W@        �       �                   �1@����X�?
             ,@        ������������������������       �                      @        �       �                     @�q�q�?             (@        ������������������������       �                     @        �       �                   �2@      �?              @        �       �                 ��Y @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 `�8"@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                   �)@���(\��?4             T@       �       �                    �?h㱪��?(            �K@        ������������������������       �                      @        �       �                 �|Y=@�&=�w��?'            �J@        �       �                   �:@�����?             5@       ������������������������       �        
             ,@        �       �                   �;@����X�?             @        ������������������������       �                     �?        �       �                   �<@r�q��?             @        ������������������������       �                     @        �       �                    $@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @@        �       �                 �|�=@ �o_��?             9@        �       �                 �|Y;@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                    @@z�G�z�?	             4@        ������������������������       �                     @        �       �                   �A@������?             .@        ������������������������       �                      @        �       �                   @D@8�Z$���?             *@        ������������������������       �                     @        �       �                    G@�q�q�?             @        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�h����?"             L@        �       �                    �?�8��8��?             (@       ������������������������       �                     $@        �       �                  �v6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     F@        �       �                    �?     ��?              H@        �       �                    �?���y4F�?             3@       �       �                 ��";@�<ݚ�?             2@        ������������������������       �                     �?        �       �                 �|�;@@�0�!��?
             1@        ������������������������       �                     �?        �       �                 `f�A@      �?	             0@       �       �                  �>@z�G�z�?             $@       �       �                 X�lE@�����H�?             "@       �       �                 �ܵ<@؇���X�?             @        ������������������������       �                     @        �       �                 ��2>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �>@����"�?             =@        �       �                   �L@�θ�?
             *@       �       �                 �|�?@r�q��?	             (@       �       �                   @>@�q�q�?             @       �       �                 `fF<@���Q��?             @        �       �                 �|�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�<@      �?
             0@        �       �                 `f�D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                 �y�/@�J�4�?             9@        �       �                  S�-@      �?              @        ������������������������       �                      @        �       �                 X�lA@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             1@        ������������������������       �                     "@        �       �                   �1@�F�j��?!            �J@        ������������������������       �                     @        �       �                 03�M@�[�IJ�?            �G@        �       �                 �|Y>@     ��?	             0@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    ;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                      @ףp=
�?             $@       �       �                   �H@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �                       @�:x@¦	^_�?             ?@       �       �                    6@������?             >@        ������������������������       �                     @        �                       `f�e@`�Q��?             9@       �       �                   �7@��.k���?             1@        ������������������������       �                     @        �       
                   �?X�Cc�?             ,@                                 �?X�<ݚ�?             "@                                 �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                 �?���Q��?             @                                 E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              	                  �G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������G�+J>�?r%�k���?[��Z���?��Z��Z�?j�a�/�?�	��7��?wwwwww�?""""""�?w�qGܱ?qG�w��?              �?�������?ZZZZZZ�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?      �?                      �?      �?                      �?�?�������?�������?333333�?t�E]t�?]t�E�?      �?      �?      �?        333333�?�������?              �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?��v`��?�Q�g���?���Q��?R���Q�?��Zk���?��RJ)��?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?      �?      �?�������?�������?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?              �?      �?        (�����?�5��P�?      �?                      �?(�����?�5��P�?              �?UUUUUU�?�������?              �?      �?      �?              �?      �?      �?              �?      �?        {	�%���?	�%����?�q�q�?r�q��?UUUUUU�?�������?�q�q�?��8��8�?              �?      �?      �?      �?                      �?              �?=��<���?�a�a�?              �?ffffff�?�������?      �?        �������?�������?      �?      �?      �?                      �?      �?        �q�q�?�q�q�?      �?        �������?�������?      �?                      �?�cj`?���8+�?              �?      �?        AZ��@�?���o)��?:����?���=��?�������?�����Ң?     ��?      �?;�;��?;�;��?      �?        �m۶m��?�$I�$I�?              �?      �?        �aܯK*�?��s���?      �?        GX�i���?�{a���?      �?        S{����?��O���?      �?        �E]t��?t�E]t�?UUUUUU�?UUUUUU�?              �?      �?        p>�cp�?������?      �?        ��+��+�?�A�A�?�Kh/��?h/�����?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?              �?      �?              �?              �?        '���?��com�?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?              �?      �?                      �?��n���?ˡE����?333333�?�������?              �?      �?        �?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?˷|˷|�?� � �?O贁N�?ƒ_,���?\���(\�?���(\��?�P^Cy�?Cy�5��?�������?UUUUUU�?� &W��?G}g����?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?        ffffff�?�����̼?־a���?��)A��?      �?        tHM0���?�x+�R�?=��<���?�a�a�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        
ףp=
�?�Q����?�������?333333�?      �?                      �?�������?�������?      �?        wwwwww�?�?              �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?              �?      �?6��P^C�?(������?9��8���?�q�q�?              �?ZZZZZZ�?�������?              �?      �?      �?�������?�������?�q�q�?�q�q�?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?                      �?      �?              �?        	�=����?�i��F�?�؉�؉�?ى�؉��?UUUUUU�?�������?UUUUUU�?UUUUUU�?�������?333333�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?              �?      �?      �?      �?              �?      �?              �?        �z�G��?{�G�z�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ��sHM�?:�&oe�?              �?���
b�?m�w6�;�?      �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?        �������?�������?�$I�$I�?۶m۶m�?              �?      �?                      �?��Zk���?�RJ)���?wwwwww�?�?      �?        ��(\���?{�G�z�?�������?�?              �?%I�$I��?�m۶m��?�q�q�?r�q��?      �?      �?      �?                      �?333333�?�������?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���bhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       n                     @v�_���?�           8�@               	                   �1@�rR���?�            �r@                                   �?XB���?             =@                                   �?      �?              @                                  �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        
       U                  x#J@�¤�h��?�             q@              L                   �K@�+2�o��?z            @h@                                  �?��l�\��?m             e@                                   �?HP�s��?!             I@                                   �?r�q��?             @                                hލC@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  �;@t��ճC�?             F@                                  �7@�<ݚ�?             "@                                  �/@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                  @E@��?^�k�?            �A@       ������������������������       �                     5@                                  @F@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@               9                     �?p�5�9��?L            �]@               8                    �?�b��[��?             �K@               7                   �G@H(���o�?            �J@       !       .                    �?~���L0�?            �H@        "       -                 `f�A@��S���?	             .@       #       ,                   @@@�q�q�?             (@       $       +                 �|�=@X�<ݚ�?             "@       %       &                 �|�;@և���X�?             @        ������������������������       �                     �?        '       *                 ��2>@      �?             @       (       )                 �ܵ<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        /       6                   �>@������?             A@       0       1                   �9@D�n�3�?             3@        ������������������������       �                     @        2       5                   �F@�q�q�?             (@       3       4                    D@z�G�z�?             $@       ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �        	             .@        ������������������������       �                     @        ������������������������       �                      @        :       ;                    �?      �?,             P@        ������������������������       �                     @        <       C                 �|�=@l�b�G��?'            �L@        =       >                   �'@��2(&�?             6@        ������������������������       �                     $@        ?       B                    �?      �?             (@       @       A                 �|�<@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        D       K                    1@��?^�k�?            �A@       E       F                   @D@�}�+r��?             3@       ������������������������       �        	             (@        G       H                 `f�)@؇���X�?             @        ������������������������       �                      @        I       J                   �F@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             0@        M       N                 `fF:@HP�s��?             9@        ������������������������       �                     $@        O       P                    �?�r����?             .@        ������������������������       �                     @        Q       T                 `f>@�<ݚ�?             "@       R       S                    N@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        V       g                 ���^@�	j*D�?5            �S@       W       f                 pf�Z@��7��?'            �N@       X       Y                    �?l��
I��?$             K@       ������������������������       �                     =@        Z       ]                    �?��H�}�?             9@        [       \                   �H@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ^       e                     �?���y4F�?             3@       _       d                   �E@      �?
             0@        `       a                 `�iJ@�q�q�?             @        ������������������������       �                      @        b       c                 03�S@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     @        h       i                    �?�IєX�?             1@       ������������������������       �        
             (@        j       m                 p�w@z�G�z�?             @        k       l                 �̒f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        o       �                    �?��P���?           �y@        p       �                 �|�=@������?N            @]@       q       �                   �8@���o� �?C            �Y@        r       y                 P��+@և���X�?             <@       s       t                    �?@4և���?
             ,@       ������������������������       �                     "@        u       v                 ���@z�G�z�?             @        ������������������������       �                      @        w       x                 ��}@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        z       }                    @d}h���?	             ,@        {       |                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ~       �                    �?�C��2(�?             &@               �                    �?r�q��?             @       �       �                     @z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��H�}�?0            �R@        �       �                 ���@�+e�X�?             9@        �       �                 �Y�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?"pc�
�?             6@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�X�<ݺ?             2@       ������������������������       �                     1@        ������������������������       �                     �?        �       �                 ���@�J�4�?             I@        ������������������������       �                     @        �       �                    �?&^�)b�?            �E@       �       �                    �?r�q��?             E@        �       �                   �<@؇���X�?             5@        ������������������������       �                     @        �       �                 �|Y=@@�0�!��?             1@        ������������������������       �                     �?        �       �                    �?      �?             0@       �       �                   @@؇���X�?             ,@        ������������������������       ����Q��?             @        ������������������������       �                     "@        ������������������������       �                      @        �       �                    �?��s����?             5@       �       �                    �?R���Q�?             4@       �       �                 �|Y=@     ��?
             0@        �       �                    ;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���@�8��8��?             (@        ������������������������       �                     @        ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                    �?����#=�?�            Pr@       �       �                 @3�.@�LQ�1	�?�            �l@       �       �                    �?���2j��?�            �i@        �       �                   �6@�q�q�?             8@        �       �                   �3@�q�q�?             (@        �       �                 P��@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?              @       �       �                 �̜!@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        �       �                 �|Y=@�8��8��?r            �f@       �       �                    �?d۬����?;            @W@       �       �                   �:@�ݜ�?3            �S@       �       �                 @3�@t�e�í�?,            �P@       �       �                 ���@ qP��B�?            �E@        �       �                 ���@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �B@        �       �                 ��Y @r�q��?             8@        �       �                   �3@���Q��?             $@        �       �                   �2@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �        
             ,@        �       �                   �;@�eP*L��?             &@        ������������������������       �                     @        �       �                 �̌!@      �?              @       ������������������������       �                     @        �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    5@��S�ۿ?             .@        �       �                 �Y�@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?`��F:u�?7            �U@       �       �                   �>@ �#�Ѵ�?6            �U@        �       �                 �|�=@����?�?            �F@       �       �                  sW@ qP��B�?            �E@        �       �                 ��,@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     C@        ������������������������       �                      @        �       �                 �?�@��p\�?            �D@       ������������������������       �                     ;@        �       �                   �?@d}h���?             ,@        ������������������������       �                      @        �       �                 @3�@�8��8��?
             (@        �       �                   �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?�	j*D�?             :@        �       �                 �|�;@��
ц��?             *@        ������������������������       �                     @        �       �                     @�q�q�?             "@       �       �                 �|Y>@      �?              @        ������������������������       �                     @        �       �                 03�1@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?8�Z$���?             *@        �       �                 �|�>@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �                          #@�b��-8�?'            �O@        �       �                 @3�4@|��?���?             ;@        ������������������������       �                     &@        �       �                    @      �?
             0@        ������������������������       �                     @                                  @�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @                                �1@�����H�?             B@                                 �?d}h���?             ,@        ������������������������       �                     @                                �0@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        	                      �̌4@���7�?             6@        
                         �?؇���X�?             @                                �=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             .@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������ *�3�?���M���?�ǉ��w�?�4
D�?�{a���?GX�i���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?KKKKKK�?iiiiii�?d���I�?7˓�4l�?��WV��?ƵHPS!�?{�G�z�?q=
ףp�?UUUUUU�?�������?      �?      �?      �?                      �?              �?t�E]t�?�E]t��?�q�q�?9��8���?      �?      �?              �?      �?                      �?�A�A�?_�_��?              �?�$I�$I�?n۶m۶�?      �?                      �?�����?�O��O��?� O	��?־a��?M0��>��?e�Cj���?����>4�?������?�?�������?�������?�������?r�q��?�q�q�?۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?      �?                      �?      �?              �?                      �?      �?        xxxxxx�?�?l(�����?(������?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?�������?333333�?      �?              �?                      �?      �?              �?      �?      �?        �Gp��?p�}��?��.���?t�E]t�?      �?              �?      �?F]t�E�?t�E]t�?      �?                      �?      �?        _�_��?�A�A�?�5��P�?(�����?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?              �?        q=
ףp�?{�G�z�?      �?        �������?�?      �?        9��8���?�q�q�?      �?      �?              �?      �?              �?        ;�;��?vb'vb'�?�y��!�?&C��6��?h/�����?Lh/����?              �?{�G�z�?
ףp=
�?UUUUUU�?�������?              �?      �?        6��P^C�?(������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?              �?        �?�?              �?�������?�������?      �?      �?              �?      �?                      �?������?�����?�C=�C=�?Xx�Wx��?r^�	��?C���?۶m۶m�?�$I�$I�?�$I�$I�?n۶m۶�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?        ]t�E�?F]t�E�?�������?UUUUUU�?�������?�������?      �?                      �?      �?              �?        {�G�z�?
ףp=
�?���Q��?R���Q�?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?/�袋.�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �q�q�?��8��8�?              �?      �?        �z�G��?{�G�z�?      �?        ���/��?�}A_��?�������?UUUUUU�?۶m۶m�?�$I�$I�?      �?        ZZZZZZ�?�������?              �?      �?      �?۶m۶m�?�$I�$I�?333333�?�������?      �?              �?        z��y���?�a�a�?333333�?333333�?      �?      �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?              �?      �?        L5����?��*�L��?��Moz��?Y�B��?�������?�������?�������?�������?�������?�������?      �?      �?              �?      �?      �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?7�p�7�?Hy�G�?\��[���?�i�i�?�1����?�rv��?��}A�?�}A_З?�������?UUUUUU�?      �?                      �?      �?        �������?UUUUUU�?333333�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?              �?        t�E]t�?]t�E�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�?�������?UUUUUU�?      �?                      �?      �?        �u�7[��?Ȥx�L��?�/����?�}A_Ч?��I��I�?l�l��?��}A�?�}A_З?�������?�������?      �?                      �?      �?              �?        �]�ڕ��?��+Q��?      �?        I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?        vb'vb'�?;�;��?�;�;�?�؉�؉�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?333333�?�������?              �?      �?                      �?;�;��?;�;��?333333�?�������?      �?                      �?      �?        �u]�u]�?QEQE�?{	�%���?	�%����?              �?      �?      �?      �?        9��8���?�q�q�?              �?      �?        �q�q�?�q�q�?I�$I�$�?۶m۶m�?      �?        F]t�E�?t�E]t�?      �?                      �?�.�袋�?F]t�E�?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ+�MhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������                           /@�s�ˈ.�?�           8�@                                   �?Ɣ��Hr�?)            �M@                                   @�G�z�?             D@        ������������������������       �                     @               
                    @h+�v:�?             A@              	                    �?      �?             8@                                @3/@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             2@        ������������������������       �        	             $@                                03�;@�\��N��?             3@        ������������������������       �                     @                                �Q��?�θ�?
             *@        ������������������������       �                      @                                    @�C��2(�?	             &@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@               d                    �?X�W9�?�           `�@               S                 pVAH@�	7���?t            `g@              &                 ���@�q�q�?Q            �_@               %                    �?��hJ,�?             A@                                 �6@6YE�t�?            �@@                                ��y@      �?              @        ������������������������       �                     @        ������������������������       �                     @               $                 �|�=@HP�s��?             9@              #                 ���@�t����?             1@              "                    �?�<ݚ�?             "@               !                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        '       8                     @�+Fi��?>             W@        (       7                    �?�q�q�?             ;@       )       ,                    �?      �?             8@        *       +                     �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        -       6                     �?R���Q�?             4@        .       /                 `f&;@�q�q�?             "@        ������������������������       �                     �?        0       5                    H@      �?              @        1       2                 �|�=@�q�q�?             @        ������������������������       �                     �?        3       4                   �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        9       @                    �?^��>�b�?+            @P@        :       ?                 X�,A@���B���?             :@       ;       <                 �|Y=@      �?             8@        ������������������������       �                     @        =       >                    �?R���Q�?
             4@       ������������������������       �        	             1@        ������������������������       �                     @        ������������������������       �                      @        A       J                    �?:�&���?            �C@        B       G                 03�-@X�Cc�?	             ,@       C       F                 �|Y=@z�G�z�?             $@        D       E                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        H       I                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        K       R                 ��(@HP�s��?             9@       L       M                 ���@�����H�?             2@        ������������������������       �                     @        N       Q                 X��A@�r����?             .@       O       P                    �?r�q��?	             (@       ������������������������       ��<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        T       U                    �?ҐϿ<��?#            �N@       ������������������������       �                     @@        V       c                    �?�c�Α�?             =@       W       Z                  �}S@����X�?             <@        X       Y                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        [       `                    �?�㙢�c�?
             7@       \       ]                 X�l@@�X�<ݺ?             2@       ������������������������       �                     (@        ^       _                 @�ys@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        a       b                 �\@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        e       �                     @�E^Y�?)           }@        f       �                    ,@h��b#��?�            �h@        g       h                   �1@p�}�ޤ�?.            @R@        ������������������������       �                      @        i       �                    �?v���EO�?-            �Q@       j       o                 `f�)@��<b���?,            @Q@       k       n                    �?�ݜ�?            �C@        l       m                   �J@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @@        p       �                   �*@�q�q�?             >@       q       x                    �?$��m��?             :@        r       s                    :@����X�?             @        ������������������������       �                     �?        t       u                    B@r�q��?             @       ������������������������       �                     @        v       w                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        y       z                 �|Y<@���y4F�?             3@        ������������������������       �                     @        {       |                 �|�=@�	j*D�?             *@        ������������������������       �                      @        }       ~                   @D@"pc�
�?             &@        ������������������������       �                     @               �                   �F@�q�q�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ��gS@������?V            �_@       �       �                    �?F�h��?E            �X@        �       �                    :@�7��?            �C@        �       �                   �E@�����H�?             2@       ������������������������       �                     "@        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        �       �                   �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        �       �                     �?6�iL�?)            �M@       �       �                    �?�L�lRT�?            �F@       �       �                    �?<=�,S��?            �A@       �       �                 ��yC@     ��?             @@       �       �                 �|�?@8�A�0��?             6@        �       �                   �@@�q�q�?             "@       �       �                   �<@      �?              @        ������������������������       �                     �?        �       �                 �|Y=@؇���X�?             @        ������������������������       �                     �?        �       �                 `fF<@r�q��?             @        ������������������������       �                     @        �       �                   �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    D@�θ�?	             *@        ������������������������       �                      @        �       �                   �Q@���!pc�?             &@       �       �                   @L@�q�q�?             "@       �       �                 ��:@      �?              @        ������������������������       �                     �?        �       �                    H@؇���X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        �       �                   �C@�z�G��?             $@        ������������������������       �                     @        �       �                    F@և���X�?             @        �       �                  x#J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        �       �                    �?@4և���?             <@       ������������������������       �                     9@        �       �                 ��n^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��F���?�            �p@        �       �                    �?���|���?%            �P@       �       �                    @���3L�?             K@       �       �                   �D@
;&����?             G@       �       �                 pf�@      �?             F@        �       �                 �|Y:@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�s��:��?             C@       �       �                 @33"@�����?             3@       �       �                 @3�@��
ц��?             *@        �       �                 pff@����X�?             @        �       �                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �8@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y>@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?D�n�3�?             3@       �       �                 �|�;@��
ц��?             *@       �       �                    4@؇���X�?             @        �       �                 �y�)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    >@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���A@      �?              @        �       �                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���0@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 ��) @P���Q�?�             i@       �       �                    �?�\=lf�?T            �`@       �       �                   @8@������?O            �_@        �       �                 ���@`���i��?             F@        �       �                 ���@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �A@        ������������������������       �        4            �T@        �       �                    3@      �?              @        ������������������������       �                     @        �       �                    5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 0SE @<���D�?,            �P@        ������������������������       �                     �?        �                          �? ����?+            @P@       �       �                    8@؇���X�?             �H@        ������������������������       �                     2@        �       �                   �;@��a�n`�?             ?@        ������������������������       �                     @        �       �                   �<@�����H�?             ;@        ������������������������       �                     "@        �                         @@@r�q��?             2@       �       �                 ���"@�q�q�?             "@        ������������������������       �                     @        �                       �|�=@���Q��?             @                                 (@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     0@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub��������������0Ȍ��?��o��?#h8����?��c+���?�������?�������?              �?xxxxxx�?�������?      �?      �?      �?      �?              �?      �?                      �?      �?        y�5���?�5��P�?              �?ى�؉��?�؉�؉�?              �?]t�E�?F]t�E�?      �?      �?              �?      �?              �?        y�%�6�?����?���=���?�ʄm�?UUUUUU�?UUUUUU�?KKKKKK�?�������?'�l��&�?e�M6�d�?      �?      �?      �?                      �?q=
ףp�?{�G�z�?<<<<<<�?�?9��8���?�q�q�?      �?      �?              �?      �?              �?              �?              �?              �?        ���,d!�?����7��?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?                      �?333333�?333333�?UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?                      �?r#7r#7�?�����?ى�؉��?��؉���?      �?      �?              �?333333�?333333�?              �?      �?              �?        �A�A�?�o��o��?%I�$I��?�m۶m��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?        q=
ףp�?{�G�z�?�q�q�?�q�q�?      �?        �������?�?�������?UUUUUU�?9��8���?�q�q�?      �?              �?              �?        mާ�d�?������?              �?5�rO#,�?�{a���?�m۶m��?�$I�$I�?�������?�������?      �?                      �?�7��Mo�?d!Y�B�?��8��8�?�q�q�?      �?        �������?UUUUUU�?      �?                      �?�������?333333�?              �?      �?              �?        �v�n���?+�"�*�?q���=�?ϩ����?�z��ի�?�
*T��?              �?�
��V�?�ԓ�ۥ�?��,d!�?��Moz��?\��[���?�i�i�?�$I�$I�?�m۶m��?              �?      �?              �?        UUUUUU�?UUUUUU�?�N��N��?vb'vb'�?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?6��P^C�?(������?      �?        vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�}��}��?AA�?Y�Cc�?T�r
^N�?�A�A�?��[��[�?�q�q�?�q�q�?              �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?ylE�pR�?'u_[�?�I��I��?l�l��?�A�A�?X|�W|��?      �?      �?/�袋.�?颋.���?UUUUUU�?UUUUUU�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?                      �?�؉�؉�?ى�؉��?              �?t�E]t�?F]t�E�?UUUUUU�?UUUUUU�?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?              �?        ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?              �?        �$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?              �?      �?        ��9����?�d\�?]t�E]�?F]t�E�?�%���^�?&���^B�?Y�B��?�Mozӛ�?      �?      �?�������?UUUUUU�?              �?      �?        �k(���?��k(��?^Cy�5�?Q^Cy��?�؉�؉�?�;�;�?�$I�$I�?�m۶m��?      �?      �?      �?                      �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?l(�����?(������?�؉�؉�?�;�;�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?UUUUUU�?      �?                      �?      �?              �?      �?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        ffffff�?�������?"=P9���?g��1��?�������?AA�?F]t�E�?F]t�E�?�q�q�?�q�q�?      �?                      �?      �?              �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        |���?|���?              �?�ȍ�ȍ�?�����?۶m۶m�?�$I�$I�?      �?        �c�1��?�s�9��?              �?�q�q�?�q�q�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJY]hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       ^                    �?�����?�           8�@               [                 p�H@*g�yw�?�            `o@                                   @Ks��?t            �f@                                   :@�KM�]�?*            �L@                                  �?@�0�!��?             A@                                  L@d}h���?             <@                               ��Y)@8�Z$���?             :@        ������������������������       �                     "@        	                          �2@������?             1@       
                           :@"pc�
�?
             &@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   -@�����H�?             "@                                 �B@      �?              @       ������������������������       �                     @                                   D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                  �7@�q�q�?             @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     7@               Z                   @B@���� �?J             _@               3                    �?�ʹ��Q�?C            �\@       !       "                    1@4և����?"             L@        ������������������������       �                     *@        #       $                    �?�^�����?            �E@        ������������������������       �                     @        %       2                    �?      �?             D@       &       )                 �̌@��G���?            �B@       '       (                   �2@ �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        *       +                    3@��
ц��?
             *@        ������������������������       �                     @        ,       -                 `�X!@���Q��?             $@        ������������������������       �                     @        .       1                 ��&@z�G�z�?             @        /       0                   �:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        4       K                    �?�Ƀ aA�?!            �M@       5       D                    �?؀�:M�?            �B@       6       =                    �?����X�?             <@        7       <                    �?؇���X�?             ,@        8       ;                 ���,@      �?             @       9       :                   �-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        >       C                 ���1@և���X�?             ,@       ?       B                 �|Y;@���!pc�?             &@        @       A                 P�@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        E       J                 `v�6@�q�q�?             "@       F       G                    0@և���X�?             @        ������������������������       �                      @        H       I                 �a2@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        L       S                 м[8@      �?             6@        M       R                    @z�G�z�?             $@       N       O                   �"@���Q��?             @        ������������������������       �                      @        P       Q                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        T       U                    �?      �?             (@        ������������������������       �                      @        V       Y                    @�z�G��?             $@        W       X                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        \       ]                    @ >�֕�?*            �Q@       ������������������������       �        (            �P@        ������������������������       �                     @        _       �                     �?�����?.           �|@        `       �                    �?��q7L��?7            �T@       a       �                    �?ꮃG��?.            @Q@       b       c                   �;@     ��?!             H@        ������������������������       �                     @        d       m                    �?�lg����?            �E@        e       l                   @G@"pc�
�?             &@       f       k                   @@@�q�q�?             @       g       j                 �|�=@z�G�z�?             @       h       i                 ��2>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        n       �                   �>@     ��?             @@       o       v                   �B@���|���?             6@       p       u                   �@@������?             .@       q       t                 `fF<@���|���?             &@       r       s                 �|�<@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        w       �                   �Q@և���X�?             @       x       y                   @E@�q�q�?             @        ������������������������       �                     �?        z                          �K@���Q��?             @       {       ~                   �G@      �?             @       |       }                 ��:@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?�q�q�?             5@       �       �                 0�"K@p�ݯ��?             3@        ������������������������       �                      @        �       �                    �?�t����?
             1@        �       �                 �U�X@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                 03�U@և���X�?             @       �       �                    C@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?X�Cc�?	             ,@       �       �                 03/O@�z�G��?             $@        ������������������������       �                     @        �       �                 tՌs@      �?             @       �       �                  DV@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    5@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�&���j�?�            �w@       �       �                    &@�ث����?�            �q@        ������������������������       �                     @        �       �                    �? ��z��?�            �q@       �       �                   �9@|(IW �?�            �q@        �       �                 �Y�@F|/ߨ�?8            @T@        �       �                    5@�C��2(�?             &@        �       �                   �2@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?`����֜?0            �Q@        ������������������������       �                     @        �       �                 0S5 @����e��?.            �P@       �       �                 @3�@г�wY;�?             A@       ������������������������       �                     ;@        �       �                   �1@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @@        �       �                   �;@���ZӼ�?             i@        �       �                     @�eP*L��?             &@        ������������������������       �                     @        �       �                  p @      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���@4z�_�\�?z            �g@        �       �                     @����?�?!            �F@        ������������������������       �                     @        �       �                 �|�=@ ���J��?            �C@       �       �                 ���@`2U0*��?             9@        ������������������������       �                     &@        �       �                    �?@4և���?
             ,@        �       �                 �|=@      �?              @        ������������������������       �                      @        ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �                     ,@        �       �                     @�ӭ�a��?Y             b@        �       �                 `f�)@\-��p�?             =@        ������������������������       �                      @        �       �                   �*@��s����?             5@       �       �                   �F@����X�?             ,@       �       �                   @D@X�<ݚ�?             "@       �       �                   @B@r�q��?             @       �       �                    @@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @@@n�����?E            �\@       �       �                    �?�4���L�?2            �U@        �       �                 P�J@�ՙ/�?             5@       �       �                 �|Y=@     ��?             0@        ������������������������       �                     �?        ������������������������       �������?             .@        �       �                 �|Y=@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|�=@��ɉ�?'            @P@       �       �                 ��) @ "��u�?             I@       ������������������������       �                     >@        �       �                 pf� @R���Q�?	             4@        ������������������������       �                      @        �       �                 ���"@�X�<ݺ?             2@        ������������������������       �                     @        �       �                    (@�C��2(�?             &@        �       �                   �<@r�q��?             @        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���!@���Q��?             .@       �       �                 @3�@�	j*D�?	             *@       �       �                 �&B@      �?              @        ������������������������       �                     �?        �       �                   �@և���X�?             @        ������������������������       �                      @        �       �                   �?@���Q��?             @        ������������������������       �                     �?        �       �                 �?�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @C@XB���?             =@        ������������������������       �        	             0@        �       �                    �?$�q-�?
             *@        ������������������������       �                     �?        �       �                   �C@�8��8��?	             (@        �       �                 ��	0@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        �                          �?|�H���?=            �V@                                  ,@�˹�m��?             C@        ������������������������       �                     �?                                 �?@-�_ .�?            �B@       ������������������������       �                     ;@                                 �?z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @                                �:@`��}3��?#            �J@              	                   �?      �?             8@        ������������������������       �                     @        
                         )@      �?             2@                                  @ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @                                 �? 	��p�?             =@        ������������������������       �                     $@                                 @�KM�]�?             3@                                  @      �?             @        ������������������������       �                     �?                                 �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     .@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������w��	�?�3����?�Tw�V�?�*�S���?�Y]���?�rS�<��?(�����?�k(���?�������?ZZZZZZ�?۶m۶m�?I�$I�$�?;�;��?;�;��?              �?�?xxxxxx�?F]t�E�?/�袋.�?      �?      �?              �?      �?        �q�q�?�q�q�?      �?      �?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?      �?              �?      �?              �?                      �?              �?B!�B�?�{����?R�0��%�?W��m�?n۶m۶�?%I�$I��?              �?֔5eMY�?�5eMYS�?      �?              �?      �?v�)�Y7�?#�u�)��?UUUUUU�?�������?      �?                      �?�؉�؉�?�;�;�?              �?333333�?�������?      �?        �������?�������?      �?      �?      �?                      �?              �?      �?        'u_�?~ylE�p�?v�)�Y7�?E>�S��?�$I�$I�?�m۶m��?�$I�$I�?۶m۶m�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?۶m۶m�?�$I�$I�?t�E]t�?F]t�E�?333333�?�������?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?�������?�������?      �?                      �?      �?              �?      �?�������?�������?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?        ffffff�?333333�?      �?      �?      �?                      �?      �?              �?        �A�A�?��+��+�?              �?      �?        �T>��u�?���(�?��\V��?��FS���?�%~F��?s��\;�?      �?      �?              �?}A_��?�}A_��?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?              �?                      �?      �?              �?      �?F]t�E�?]t�E]�?�?wwwwww�?F]t�E�?]t�E]�?�������?�������?              �?      �?                      �?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?Cy�5��?^Cy�5�?      �?        �������?�������?�������?�������?              �?      �?        ۶m۶m�?�$I�$I�?333333�?�������?              �?      �?                      �?              �?%I�$I��?�m۶m��?ffffff�?333333�?      �?              �?      �?      �?      �?              �?      �?                      �?      �?      �?              �?      �?        %�,.�j�?k�LG�U�?fI9 2�?�ϴ5�n�?              �?ǬӢ�~�?șb��
�?�p$�Ax�?Bx�>�=�?�Hx�5�?�����H�?]t�E�?F]t�E�?      �?      �?      �?              �?      �?              �?      �?              �?        �������?�A�A�?      �?        �>����?|���?�?�?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?        \���(\�?���(\��?]t�E�?t�E]t�?      �?              �?      �?      �?                      �?����?t���G'�?��I��I�?l�l��?      �?        ��-��-�?�A�A�?���Q��?{�G�z�?      �?        n۶m۶�?�$I�$I�?      �?      �?      �?        �������?UUUUUU�?      �?              �?        �q�q�?�8��8��?a����?�{a���?      �?        z��y���?�a�a�?�m۶m��?�$I�$I�?r�q��?�q�q�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?              �?        �K*���?A�V���?kʚ����?S֔5eM�?�<��<��?�a�a�?      �?      �?              �?wwwwww�?�?�������?333333�?              �?      �?        �����?�����?�G�z�?���Q��?      �?        333333�?333333�?              �?��8��8�?�q�q�?      �?        ]t�E�?F]t�E�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        333333�?�������?vb'vb'�?;�;��?      �?      �?      �?        ۶m۶m�?�$I�$I�?              �?333333�?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?GX�i���?�{a���?      �?        �؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?              �?              �?        y��x���?�!�!�?��P^Cy�?^Cy�5�?              �?S�n0E�?к����?      �?        �������?�������?              �?      �?        �琚`��?M0��>��?      �?      �?              �?      �?      �?�������?�������?              �?      �?              �?        ������?�{a���?      �?        �k(���?(�����?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ4
hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       p                    �?��eC~�?�           8�@               '                     @����X�?�            �o@                                  @Tۢ��(�?V            �`@        ������������������������       �                     �?                                   �?t�e�í�?U            �`@                                   �? ���J��?            �C@              
                 0Cd=@�?�|�?            �B@               	                 03[:@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �@@        ������������������������       �                      @               $                    L@�¦�{��?9            �W@              #                    :@$�q-�?7            �V@              "                    �?H�ՠ&��?             K@                                 �'@؇���X�?            �H@        ������������������������       �                     .@                                  �*@H�V�e��?             A@                                   <@�q�q�?             (@        ������������������������       �                     @                                  �B@�����H�?             "@       ������������������������       �                     @                                   D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?��2(&�?             6@        ������������������������       �                     "@               !                   �E@�θ�?             *@                                   <@�C��2(�?             &@                                  �9@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �B@        %       &                     �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        (       Q                    �?�O
��?G            @]@       )       4                 �̌@b�2�tk�?+             R@        *       3                    �?�חF�P�?             ?@       +       .                 ���@д>��C�?             =@        ,       -                 �|Y:@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        /       0                    �?���7�?             6@       ������������������������       �                     4@        1       2                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        5       <                  �#@�>$�*��?            �D@        6       ;                 @3�@@4և���?             ,@        7       8                 �?�@؇���X�?             @        ������������������������       �                     �?        9       :                   �9@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        =       B                    �?��}*_��?             ;@        >       ?                   �-@և���X�?             @        ������������������������       �                      @        @       A                 ���,@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        C       D                    �?�z�G��?             4@        ������������������������       �                     @        E       L                 �|�;@���Q��?
             .@       F       G                    '@      �?              @        ������������������������       �                      @        H       K                    4@r�q��?             @       I       J                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        M       N                   �>@؇���X�?             @        ������������������������       �                     @        O       P                 ���0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        R       k                    @������?            �F@       S       Z                    �?      �?             D@        T       Y                    �?z�G�z�?             @       U       V                    �?      �?             @        ������������������������       �                      @        W       X                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        [       b                 ���4@��R[s�?            �A@        \       ]                    �?      �?              @        ������������������������       �                     @        ^       _                    -@z�G�z�?             @        ������������������������       �                     @        `       a                 `fv1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        c       f                 �̼6@�>����?             ;@        d       e                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        g       h                    @���7�?             6@       ������������������������       �                     0@        i       j                    @r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        l       o                    @���Q��?             @       m       n                   @C@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        q       �                    �?"~��F��?$           �|@       r       �                    �?X�9H���?�             w@        s       �                    �?@�0�!��?"            �I@       t       }                 �|Y<@؇���X�?             E@        u       z                 �܅6@�q�q�?             (@        v       y                 hfF&@r�q��?             @       w       x                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        {       |                  �}S@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ~                        `f�3@(;L]n�?             >@       ������������������������       �                     1@        �       �                   @@@$�q-�?	             *@        ������������������������       �                      @        �       �                   �A@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �C@�q�q�?             "@       �       �                    .@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     �?$}3���?�            �s@        �       �                 03:@�^�����?!             O@        ������������������������       �                     @        �       �                   �E@6C�z��?            �L@       �       �                    �?      �?             D@       �       �                 ��yC@�f7�z�?             =@       �       �                 �|�<@�KM�]�?             3@        ������������������������       �                      @        �       �                 �|�?@"pc�
�?             &@        �       �                   �>@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                  x#J@���!pc�?             &@        ������������������������       �                     �?        �       �                    7@z�G�z�?             $@        ������������������������       �                     �?        �       �                    A@�����H�?             "@        ������������������������       �                     @        �       �                   �B@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �G@������?
             1@        ������������������������       �                      @        �       �                   �J@X�<ݚ�?             "@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @���?�            p@        �       �                    4@�nkK�?/            @Q@        �       �                   �2@r�q��?             @        ������������������������       �                      @        �       �                   �'@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        �       �                    �?�i�y�?*            �O@       �       �                    �?@9G��?"            �H@        ������������������������       �                     �?        �       �                    F@ �q�q�?!             H@       �       �                   @D@�X�<ݺ?             B@       �       �                 �|�=@г�wY;�?             A@        �       �                   �'@      �?             0@        ������������������������       �                     "@        �       �                   �3@؇���X�?             @       �       �                 �|�<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �      �?              @        ������������������������       �        	             (@        ������������������������       �                     ,@        �       �                   �:@�D�az�?}            �g@        �       �                    �?`����֜?3            �Q@        ������������������������       �                     �?        �       �                   @4@@	tbA@�?2            @Q@        �       �                   �3@(;L]n�?             >@       ������������������������       �                     2@        �       �                    �?�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                    �C@        �       �                    �?�j��b�?J            �]@       �       �                  s�@$	4�}�?C            �Z@        ������������������������       �                     1@        �       �                 ��@�r����?8            �V@        �       �                 �|Y=@�z�G��?             $@        ������������������������       �                     �?        �       �                 X�I@�<ݚ�?             "@       ������������������������       �����X�?             @        ������������������������       �                      @        �       �                    �?���(\��?1             T@        ������������������������       �                     �?        �       �                 pf� @���!���?0            �S@       �       �                   �@�8��8��?#             N@        �       �                   @@@     ��?             0@       �       �                   �?@�z�G��?             $@       �       �                 �|�<@      �?              @        ������������������������       �                     @        �       �                 �|Y>@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �?�@���7�?             F@        ������������������������       �                     5@        �       �                 @3�@���}<S�?             7@        �       �                   �A@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     3@        �       �                    (@���y4F�?             3@       �       �                   �?@�	j*D�?             *@       �       �                 ���"@      �?              @        �       �                 0S%"@      �?             @       �       �                 �|Y<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        �                           @�μ���?5            @V@        �                          �?�q�q�?            �C@       �       �                    :@������?             >@        �       �                    �?X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        �                            �?؇���X�?             5@       �       �                   �7@d}h���?	             ,@        ������������������������       �                      @        �       �                 �̾w@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     @              	                    �?X�<ݚ�?             "@                                @      �?             @                                �?�q�q�?             @                                6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        
                         �?���Q��?             @                               �2@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                  @j�q����?             I@                                0@����X�?             <@                             ��-@�n_Y�K�?             *@                                &@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     .@                                 @���7�?             6@                                �?�8��8��?	             (@       ������������������������       �                      @                                 @      �?             @        ������������������������       �                      @                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub���������������Kkz�?�fh)�?�$I�$I�?�m۶m��?�M1j�۴?Hֹ�d�?      �?        �rv��?�1����?�A�A�?��-��-�?к����?*�Y7�"�?      �?      �?              �?      �?                      �?              �?��v�@�?�-q���?;�;��?�؉�؉�?{	�%���?������?�$I�$I�?۶m۶m�?              �?ZZZZZZ�?iiiiii�?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?t�E]t�?��.���?              �?�؉�؉�?ى�؉��?F]t�E�?]t�E�?�������?�������?              �?      �?                      �?      �?                      �?              �?      �?      �?              �?      �?        �
��
��?���?9��8���?�8��8��?��RJ)��?�Zk����?|a���?a���{�?�$I�$I�?۶m۶m�?              �?      �?        F]t�E�?�.�袋�?              �?      �?      �?              �?      �?                      �?�18���?�����?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?      �?                      �?      �?        B{	�%��?_B{	�%�?�$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?        333333�?ffffff�?              �?�������?333333�?      �?      �?              �?�������?UUUUUU�?      �?      �?              �?      �?              �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?        wwwwww�?�?      �?      �?�������?�������?      �?      �?      �?              �?      �?              �?      �?              �?        X|�W|��?PuPu�?      �?      �?              �?�������?�������?              �?      �?      �?      �?                      �?�Kh/��?h/�����?�������?�������?      �?                      �?�.�袋�?F]t�E�?      �?        �������?UUUUUU�?              �?      �?        333333�?�������?      �?      �?              �?      �?              �?        �A^%���?���j�1�?G��*iT�?�*iT[��?ZZZZZZ�?�������?۶m۶m�?�$I�$I�?�������?�������?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�?      �?        �؉�؉�?;�;��?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?                      �?
ςc|�?����q�?!�B�?���{��?      �?        ��Gp�?~��G�?      �?      �?a���{�?O#,�4��?(�����?�k(���?              �?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        t�E]t�?F]t�E�?      �?        �������?�������?      �?        �q�q�?�q�q�?              �?�������?�������?      �?                      �?xxxxxx�?�?      �?        r�q��?�q�q�?�������?�������?              �?      �?              �?        ����? ���?�Mozӛ�?d!Y�B�?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?        �������?AA�?������?9/���?      �?        �������?UUUUUU�?��8��8�?�q�q�?�?�?      �?      �?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?              �?              �?      �?      �?              �?        W�+���?G}g����?�������?�A�A�?      �?        �%~F��?ہ�v`��?�������?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �N��?��/���?��bEi�?�@�Ե�?      �?        �������?�?ffffff�?333333�?              �?9��8���?�q�q�?�m۶m��?�$I�$I�?      �?        ffffff�?�����̼?      �?        ��	�Z�?T:�g *�?UUUUUU�?UUUUUU�?      �?      �?ffffff�?333333�?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �.�袋�?F]t�E�?      �?        ӛ���7�?d!Y�B�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?        6��P^C�?(������?vb'vb'�?;�;��?      �?      �?      �?      �?      �?      �?              �?      �?              �?              �?      �?      �?                      �?      �?              �?              �?        �\��?�я~���?UUUUUU�?UUUUUU�?wwwwww�?�?�q�q�?r�q��?              �?      �?        ۶m۶m�?�$I�$I�?I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?r�q��?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        �������?333333�?      �?      �?              �?      �?              �?        =
ףp=�?
ףp=
�?�m۶m��?�$I�$I�?ى�؉��?;�;��?�m۶m��?�$I�$I�?              �?      �?                      �?      �?        �.�袋�?F]t�E�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��;hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                 �J/@���%&�?�           8�@                                 �,@������?�            @x@                                ��-@�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?               5                    �?l=.�5�?�            �w@                                ���@n>�X�q�?8             W@                                  �6@r�q��?             >@        	                           �?      �?             @       
                           5@���Q��?             @                               �{@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                0��@�8��8��?             8@                               ��Y@ףp=
�?             4@        ������������������������       �                     @                                ���@�t����?
             1@                                  �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                                �|�=@      �?              @                               �|�:@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @               &                   P,@`՟�G��?%             O@              %                 �F$*@\X��t�?             G@                                   �?�G��l��?             E@        ������������������������       �                     1@        !       "                     @z�G�z�?             9@        ������������������������       �                     @        #       $                 �|Y=@�GN�z�?             6@        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                     @        '       (                     @      �?	             0@        ������������������������       �                     �?        )       0                    �?�r����?             .@       *       /                    �?      �?              @       +       .                 ���,@�q�q�?             @       ,       -                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        1       2                    �?؇���X�?             @        ������������������������       �                     @        3       4                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        6       c                 ��) @6�����?�            �q@       7       b                    @���.n�?\            �c@       8       ]                    �?�-���?[            `c@       9       H                   �3@�L���?V            �b@        :       E                   �2@     ��?
             0@       ;       <                    �?�<ݚ�?             "@        ������������������������       �                     �?        =       @                   �0@      �?              @        >       ?                 pf�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        A       B                   �1@z�G�z�?             @        ������������������������       �                     �?        C       D                 ��@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        F       G                 �?�@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        I       J                     @�5[|/��?L            �`@        ������������������������       �                     ,@        K       N                   �7@�1e�3��?E            �]@        L       M                    �?�LQ�1	�?             7@        ������������������������       �                     @        ������������������������       �                     4@        O       \                   �@@��s��?7            �W@       P       Y                    ?@�IєX�?'             Q@       Q       R                 �|Y=@��ɉ�?%            @P@        ������������������������       �                     :@        S       X                  sW@�7��?            �C@        T       U                    �?r�q��?             (@        ������������������������       �                     �?        V       W                 ��,@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     ;@        Z       [                 P�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        ^       a                    �?����X�?             @        _       `                 P�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        d       �                    �?l��э�?N            �_@       e       j                   �4@�"'`�]�?E            @\@        f       i                    �?HP�s��?             9@       g       h                    �? �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                     �?        k       �                   @@@      �?6             V@       l       �                 �|�=@��.k���?!            �I@       m       �                    �?�ʻ����?             A@       n       o                   �5@     ��?             @@        ������������������������       �                      @        p       s                    �?d��0u��?             >@        q       r                     @���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        t       u                 @3"@`�Q��?             9@        ������������������������       �                     @        v       w                   �<@��s����?             5@       ������������������������       �                      @        x       {                     @�	j*D�?             *@        y       z                   �'@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        |                           (@�����H�?             "@        }       ~                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�t����?	             1@        ������������������������       �                     $@        �       �                     @����X�?             @       ������������������������       �                     @        �       �                 ���!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�MI8d�?            �B@        �       �                 `f�&@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     >@        ������������������������       �        	             ,@        �       �                    �?�� ���?�            0t@        �       �                    @tk~X��?]             b@       �       �                 0#
9@�N̸��?R            �_@        �       �                    �?������?             ;@       �       �                    �?"pc�
�?             6@        �       �                     @X�<ݚ�?             "@       �       �                   �6@����X�?             @       �       �                   �2@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        �       �                 X��D@���Q��?             @       �       �                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @ "��u�?B             Y@       �       �                    �?@��8��?>             X@       ������������������������       �        5            @T@        �       �                    �?�r����?	             .@        ������������������������       �                      @        �       �                    @8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        �       �                    @�t����?             1@       �       �                    �?"pc�
�?             &@        ������������������������       �                     @        �       �                 ��T?@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �                       ��!T@��Ж�H�?l            `f@       �       �                     �?�G�z��?`             d@        �       �                  �>@�)��V��?0            �T@        �       �                    �?�q�q�?             >@       �       �                 ��$:@8^s]e�?             =@        ������������������������       �                      @        �       �                    �?������?             ;@        �       �                 ��";@      �?             (@        ������������������������       �                      @        �       �                 �ܵ<@�z�G��?             $@        ������������������������       �                     �?        �       �                 ���=@�<ݚ�?             "@       �       �                 X��E@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �Q@������?	             .@       �       �                   @>@�q�q�?             (@       �       �                 `fF<@���Q��?             $@       �       �                 03k:@�q�q�?             "@        ������������������������       �                     �?        �       �                   �K@      �?              @       �       �                    H@����X�?             @       �       �                 �|�<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 0�"K@�c�����?            �J@       �       �                    �?     ��?             @@        �       �                 p�i@@և���X�?             @        �       �                  �>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�<@HP�s��?             9@        �       �                    7@���Q��?             @        ������������������������       �                      @        �       �                   �;@�q�q�?             @        ������������������������       �                     �?        �       �                 `f�D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        �       �                    �?�ՙ/�?             5@       �       �                   �L@�eP*L��?             &@       �       �                   �8@�q�q�?             "@        �       �                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @C@z�G�z�?             $@        �       �                    >@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �                          @"pc�
�?0            @S@       �       �                    �?����|e�?%             K@       �       �                     @H%u��?             9@        ������������������������       �                     "@        �       �                 �|�>@     ��?             0@       �       �                 �|=@$�q-�?	             *@       ������������������������       �                      @        �       �                 м�5@z�G�z�?             @        ������������������������       �                     @        �       �                 0��C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �T)D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �                           )@J�8���?             =@        ������������������������       �                     "@                                 �?P���Q�?             4@                             8#�1@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     $@                                 �?�nkK�?             7@        ������������������������       �                     $@                              pf�C@$�q-�?             *@        	      
                   @z�G�z�?             @        ������������������������       �                      @                                 @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                �H@p�ݯ��?             3@                                :@؇���X�?	             ,@        ������������������������       �                     @                                 �?����X�?             @                                �?���Q��?             @                                �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������g *��?�0���M�?���:*�??��W�?UUUUUU�?UUUUUU�?              �?      �?        ���Q���?r1����?�B����?ozӛ���?�������?UUUUUU�?      �?      �?333333�?�������?      �?      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?�������?�������?      �?        <<<<<<�?�?�q�q�?�q�q�?              �?      �?              �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?        �1�c��?�s�9��?��Moz��?!Y�B�?��y��y�?1�0��?              �?�������?�������?      �?        �袋.��?]t�E�?              �?      �?                      �?      �?      �?      �?        �������?�?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        H���@�?��.�d��?��Ѐ%��?Kz���?=���?�qa�?}���g�?L�Ϻ��?      �?      �?9��8���?�q�q�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?              �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?                      �?N6�d�M�?'�l��&�?      �?        �/���?W'u_�?��Moz��?Y�B��?              �?      �?        q�����?�X�0Ҏ�?�?�??�?��? �����?      �?        ��[��[�?�A�A�?�������?UUUUUU�?      �?        /�袋.�?F]t�E�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?��r�\.�?i4�F��?zja���?+=����?q=
ףp�?{�G�z�?�������?UUUUUU�?              �?      �?                      �?      �?      �?�?�������?�������?<<<<<<�?      �?      �?              �?DDDDDD�?wwwwww�?�������?333333�?              �?      �?        ��(\���?{�G�z�?              �?z��y���?�a�a�?      �?        vb'vb'�?;�;��?      �?      �?      �?                      �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?                      �?�������?�������?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?��L���?L�Ϻ��?�$I�$I�?۶m۶m�?      �?                      �?      �?              �?        a�E8S�?�~ �cV�?9��8���?r�q��?�F��h4�?.���r��?{	�%���?B{	�%��?F]t�E�?/�袋.�?�q�q�?r�q��?�$I�$I�?�m۶m��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?333333�?�������?      �?      �?      �?                      �?              �?���Q��?�G�z�?UUUUUU�?UUUUUU�?              �?�?�������?              �?;�;��?;�;��?      �?                      �?      �?        <<<<<<�?�?/�袋.�?F]t�E�?      �?              �?      �?      �?                      �?      �?        J���s�?k��P�?�������?�������?]V��F�?GS��r�?UUUUUU�?UUUUUU�?	�=����?|a���?      �?        {	�%���?B{	�%��?      �?      �?              �?333333�?ffffff�?      �?        �q�q�?9��8���?�$I�$I�?�m۶m��?              �?      �?                      �?�?wwwwww�?UUUUUU�?UUUUUU�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?              �?                      �?              �?      �?        �V�9�&�?:�&oe�?      �?      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?        q=
ףp�?{�G�z�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        �<��<��?�a�a�?]t�E�?t�E]t�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        �������?�������?      �?      �?      �?                      �?      �?        /�袋.�?F]t�E�?����K�?	�%����?)\���(�?���Q��?      �?              �?      �?�؉�؉�?;�;��?      �?        �������?�������?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�rO#,��?|a���?              �?ffffff�?�������?�������?�������?              �?      �?              �?        �Mozӛ�?d!Y�B�?      �?        �؉�؉�?;�;��?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        Cy�5��?^Cy�5�?�$I�$I�?۶m۶m�?              �?�$I�$I�?�m۶m��?�������?333333�?      �?      �?              �?      �?              �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJS�)/hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                    �?�Wa�O�?�           8�@              K                     @*���M��?5           �}@                                  �1@���E��?�            �k@        ������������������������       �        	             .@               >                 ��UO@��>��?            �i@              7                   �J@>��"��?f            �e@                                  �?:%�[��?U            �a@                                   �?������?            �D@       	       
                   �B@ >�֕�?            �A@       ������������������������       �                     :@                                0#R;@�<ݚ�?             "@                                 �'@      �?              @        ������������������������       �                     @                                    �?      �?             @        ������������������������       �                      @                                  �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               4                   �G@0�W���?;            @Y@                               `fF:@�A����?7             W@       ������������������������       �        "            �L@               +                  Y>@">�֕�?            �A@              "                 ��";@     ��?             0@                               �|�<@�q�q�?             "@        ������������������������       �                      @                                �|�?@և���X�?             @        ������������������������       �                      @                                   �?z�G�z�?             @        ������������������������       �                     �?                !                   �C@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        #       $                   �;@և���X�?             @        ������������������������       �                      @        %       &                 �|Y=@z�G�z�?             @        ������������������������       �                      @        '       *                 X��B@�q�q�?             @       (       )                 0C�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ,       3                   �B@�KM�]�?
             3@        -       2                   �A@      �?              @       .       1                    �?؇���X�?             @       /       0                  �>@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        5       6                 `f�3@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        8       ;                    �?��� ��?             ?@        9       :                   �L@      �?             @        ������������������������       �                      @        ������������������������       �                      @        <       =                   �R@�>����?             ;@       ������������������������       �                     9@        ������������������������       �                      @        ?       D                 `fmj@���!pc�?            �@@       @       A                    �?�LQ�1	�?             7@       ������������������������       �                     3@        B       C                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        E       H                    �?���Q��?             $@        F       G                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        I       J                   �?@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        L       o                    �? ���m>�?�            p@        M       \                 �̌@���H.�?#             I@       N       U                    �?r�q��?             8@       O       T                    �?�t����?             1@       P       S                 ���@      �?             0@        Q       R                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?        V       W                 ���@����X�?             @        ������������������������       �                     @        X       Y                   �9@�q�q�?             @        ������������������������       �                     �?        Z       [                 �Y5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ]       f                 ��&@$��m��?             :@        ^       e                    �?8�Z$���?             *@       _       `                    9@�8��8��?             (@       ������������������������       �                      @        a       d                 03�!@      �?             @       b       c                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        g       n                    @��
ц��?	             *@       h       i                    �?�z�G��?             $@        ������������������������       �                     @        j       m                    �?և���X�?             @       k       l                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        p       q                    $@�_�/�?�            �i@        ������������������������       �                      @        r       �                   �C@���x��?�            �i@       s       �                 ��q1@�I�,ѽ�?|            @g@       t       �                    �?@�qmNh�?w            `f@        u       v                   �6@�GN�z�?             6@        ������������������������       �                     @        w       x                 ���@�KM�]�?             3@        ������������������������       �                     "@        y       �                 �|�=@z�G�z�?             $@       z       }                   @@����X�?             @       {       |                 �|=@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ~                        �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���@P��-�?i            �c@        ������������������������       �                     1@        �       �                   @C@ �Cc}�?^            �a@       �       �                    �?�:�^���?\            �`@        �       �                 �|Y=@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        �       �                 ���@85�}C�?T            �^@        ������������������������       �                     @        �       �                 �?�@�IєX�?S            �]@        �       �                   �@�]0��<�?)            �N@       �       �                 P�N@�IєX�?             A@       �       �                 �|�<@XB���?             =@       ������������������������       �                     3@        �       �                 �|Y>@ףp=
�?             $@       �       �                 pf�@      �?              @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                    >@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ;@        �       �                 0SE @��ϭ�*�?*             M@        �       �                 ��) @؇���X�?             <@       �       �                 @3�@$�q-�?             :@        �       �                    :@z�G�z�?             @        ������������������������       �                      @        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �4@���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                      @        �       �                 �|�=@(;L]n�?             >@       ������������������������       �                     ;@        �       �                 ��)"@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       ����Q��?             @        �       �                 �|�;@և���X�?             @       �       �                    �?      �?             @       �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        �       �                    �?��C:��?�             m@       �       �                     @�z�G��?J             ^@       �       �                 03�a@ >�֕�?*            �Q@       �       �                    �?�]0��<�?$            �N@       �       �                    �?���U�?"            �L@        ������������������������       �                     7@        �       �                    �?�IєX�?             A@        �       �                   �7@�t����?
             1@        ������������������������       �                     �?        �       �                     �?      �?	             0@        ������������������������       �                     @        �       �                   �E@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     @        �       �                    $@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                    @��H�}�?              I@       �       �                    @��Zy�?            �C@        ������������������������       �                     @        �       �                    �?ҳ�wY;�?             A@        �       �                    �?z�G�z�?             $@       �       �                    �?      �?              @        �       �                    �?���Q��?             @       �       �                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?r�q��?             8@        �       �                    @@�q�q�?             "@       �       �                    �?      �?              @       �       �                    4@����X�?             @        ������������������������       �                     �?        �       �                 �|�;@r�q��?             @        ������������������������       �                     @        �       �                 ��1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��T?@��S�ۿ?             .@       ������������������������       �                      @        �       �                   �7@؇���X�?             @        ������������������������       �                     @        �       �                   �E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @�C��2(�?             &@        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    @��o���?I            @\@        �       �                     @������?             .@        ������������������������       �                     @        �       �                     @      �?              @        ������������������������       �                     @        �       �                    @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          G@�[$�G�?>            �X@       �                          @�k��?7            @V@       �                       �|�=@z���=��?.            @S@       �       �                     �?r�qG�?             H@        �       �                    �?�q�q�?             (@        �       �                 �U�X@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    7@և���X�?             @        ������������������������       �                      @        �       �                 ���M@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                                  )@r�q��?             B@        ������������������������       �                     �?                               �v6@؇���X�?            �A@             
                ��.@HP�s��?             9@                               �4@�r����?             .@                              P�@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?              	                03�-@�8��8��?
             (@       ������������������������       �        	             &@        ������������������������       �                     �?        ������������������������       �                     $@                              03�7@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     =@        ������������������������       �        	             (@                                �H@�q�q�?             "@        ������������������������       �                     @                                 �?      �?             @        ������������������������       �                     �?                                �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������M}<���?g�/��?1N�����?�c�D@|�?�G��G��?]p�\p��?              �?�	����?����?�����?��R�O2�?+l$Za�?�'�K=�?������?p>�cp�?�A�A�?��+��+�?              �?�q�q�?9��8���?      �?      �?              �?      �?      �?              �?      �?      �?      �?                      �?      �?                      �?�&��?���g��?C���,�?�Mozӛ�?      �?        _�_��?�A�A�?      �?      �?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?      �?              �?      �?      �?�$I�$I�?۶m۶m�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �k(���?(�����?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�{����?�B!��?      �?      �?      �?                      �?�Kh/��?h/�����?      �?                      �?t�E]t�?F]t�E�?Y�B��?��Moz��?              �?      �?      �?              �?      �?        333333�?�������?      �?      �?              �?      �?        �������?UUUUUU�?      �?                      �?�F�F�F�?����?�z�G��?���(\��?UUUUUU�?�������?�?<<<<<<�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�N��N��?vb'vb'�?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?              �?      �?              �?                      �?�؉�؉�?�;�;�?333333�?ffffff�?              �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?      �?        m��Š"�?�<���?              �?i\���h�?���Ѹ�?,���?��~�駿?I=W�l�?�Fu��?�袋.��?]t�E�?              �?�k(���?(�����?      �?        �������?�������?�m۶m��?�$I�$I�?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        6��(S��?R��fu�?      �?        %I�$I��?۶m۶m�?}�'}�'�?l�l��?;�;��?;�;��?              �?      �?        �}�K�`�?������?              �?�?�?\2�h��?;ڼOqɠ?�?�?GX�i���?�{a���?      �?        �������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?      �?                      �?      �?        ����=�?|a���?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��y��y�?�a�a�?              �?      �?                      �?�������?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?�$I�$I�?۶m۶m�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?        -����W�?����4P�?333333�?ffffff�?�A�A�?��+��+�?;ڼOqɠ?\2�h��?p�}��?	�#����?              �?�?�?�?<<<<<<�?      �?              �?      �?              �?;�;��?�؉�؉�?              �?      �?                      �?              �?�q�q�?9��8���?      �?                      �?{�G�z�?
ףp=
�?� � �?\��[���?              �?�������?�������?�������?�������?      �?      �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?�?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ]t�E�?F]t�E�?      �?      �?      �?                      �?      �?         x�!��?��	���?�?wwwwww�?              �?      �?      �?              �?�������?�������?      �?                      �?s
^N���?4և����?��MmjS�?+Y�JV��?�cj`��?
qV~B��?UUUUUU�?UUUUUU�?�������?�������?�������?�������?              �?      �?        �$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?        �������?UUUUUU�?              �?۶m۶m�?�$I�$I�?q=
ףp�?{�G�z�?�������?�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ffffff�?333333�?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ[س=hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       ^                    �?H���I�?�           8�@                                    @@�j���?�            @o@                                  @Pa�	�?V            �`@        ������������������������       �                     �?                                   �?�z�N��?U            ``@                                0Cd=@`Ql�R�?             �G@               
                    �?r�q��?             @              	                 03[:@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �D@                                   �?�Ń��̧?5             U@                                   �? �q�q�?             H@        ������������������������       �                     5@                                `f&'@�>����?             ;@                                  �J@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                  �;@���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     B@               '                 �̌@�m����?M            �]@                                pff@      �?             @@                                 s@      �?             @       ������������������������       �                     @        ������������������������       �                     �?               &                   �9@h�����?             <@                                ��@�C��2(�?             &@        ������������������������       �                     @                %                    �?z�G�z�?             @       !       $                 P�N@      �?             @       "       #                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     1@        (       3                    @8�$�>�?8            �U@        )       *                    �?�<ݚ�?             "@        ������������������������       �                     @        +       ,                    �?���Q��?             @        ������������������������       �                     �?        -       0                    �?      �?             @        .       /                 @3�2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       2                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        4       5                   �-@x�(�3��?1            @S@        ������������������������       �                     "@        6       7                    /@.Lj���?,             Q@        ������������������������       �                      @        8       ]                 ��Y7@�X����?+            �P@       9       X                    �?��V�I��?            �G@       :       M                 �|Y=@�D����?             E@       ;       <                    �?���B���?             :@        ������������������������       �                      @        =       F                  �#@�q�q�?             8@       >       E                 pf� @�C��2(�?             &@        ?       D                    �?r�q��?             @       @       A                 �?�@z�G�z�?             @        ������������������������       �                     @        B       C                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        G       L                    �?�	j*D�?             *@        H       I                 �[$@�q�q�?             @        ������������������������       �                      @        J       K                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        N       W                   @B@      �?             0@       O       V                 �|�=@؇���X�?	             ,@       P       U                    �?      �?              @       Q       T                    �?����X�?             @        R       S                 P�h2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        Y       \                    @z�G�z�?             @       Z       [                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     3@        _                       �U�R@�7�&,��?           �|@       `       �                     �?��b7E�?           �{@        a       ~                   �B@z�G�z�?)            @P@       b       }                    �?������?            �D@       c       j                    �?4�B��?            �B@        d       e                    <@����X�?             @        ������������������������       �                     �?        f       g                  �>@r�q��?             @        ������������������������       �                     @        h       i                   �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        k       l                   �<@�q�q�?             >@        ������������������������       �                     @        m       |                    R@�θ�?             :@       n       {                   �K@r�q��?             8@       o       p                 �̌/@������?             1@        ������������������������       �                     @        q       z                   �>@�q�q�?	             (@       r       y                   @G@      �?              @       s       x                 X��B@�q�q�?             @       t       u                 `fF<@      �?             @        ������������������������       �                     �?        v       w                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @               �                    �? �q�q�?             8@        ������������������������       �                     &@        �       �                   �G@$�q-�?	             *@       ������������������������       �                     $@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?������?�            �w@       �       �                    ,@(32v�c�?�            `t@        �       �                    '@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    A@�q�D�?�            0t@       �       �                 �Y�@D�2y�?�            0p@        �       �                     @�<ݚ�?            �F@        ������������������������       �                      @        �       �                   �3@>��C��?            �E@        ������������������������       �                      @        �       �                   �6@����X�?            �A@        �       �                    5@�q�q�?             @        �       �                 P�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?V�a�� �?             =@       �       �                    �?�J�4�?             9@       �       �                 ���@r�q��?             8@       ������������������������       �                     $@        �       �                 �|=@����X�?             ,@        ������������������������       �                     @        ������������������������       ����Q��?             $@        ������������������������       �                     �?        �       �                    =@      �?             @       �       �                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �>@��8����?�            �j@       �       �                    �?P��a4�?u            �g@        �       �                     @�8��8��?             B@        ������������������������       �                     @        �       �                    �?ףp=
�?             >@       �       �                 03s@�LQ�1	�?             7@       �       �                 ���@�����?             5@        ������������������������       �                     @        �       �                 ��(@      �?             0@       ������������������������       �؇���X�?             ,@        ������������������������       �                      @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @�}�+r��?`             c@        �       �                 �|Y=@`Jj��?             ?@       ������������������������       �                     7@        �       �                 �|�=@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?����&!�?K            @^@       �       �                    �?�7��?H            @]@       �       �                    9@�f�¦ζ?C            �Z@        �       �                 0S5 @P����?!            �M@       �       �                   �1@Pa�	�?            �@@        ������������������������       ��q�q�?             @        ������������������������       �                     >@        ������������������������       �                     :@        �       �                   �;@�8��8��?"             H@        �       �                   �:@և���X�?             @        �       �                 �T@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �� @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y=@��Y��]�?            �D@        ������������������������       �                     "@        �       �                 �|�=@      �?             @@       �       �                  sW@�g�y��?             ?@        �       �                 pf�@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     ;@        ������������������������       �                     �?        �       �                    6@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                    �?���B���?             :@       �       �                 `fF)@�q�q�?             8@       �       �                     @�KM�]�?             3@        ������������������������       �                     @        �       �                   �?@؇���X�?
             ,@        �       �                 pff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @@@�8��8��?             (@        �       �                 P�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 0�_A@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �?�@      �?&             P@        ������������������������       �                     3@        �       �                 @3�@`Ӹ����?            �F@        ������������������������       �                     �?        �       �                   �E@`���i��?             F@        �       �                    �?�nkK�?             7@       �       �                   �)@�X�<ݺ?
             2@        ������������������������       �                     *@        �       �                     @z�G�z�?             @       �       �                   @D@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        �       �                    @      �?             J@        �       �                   �C@      �?             0@       �       �                    �?r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        �                          �?�8��8��?             B@        �                          P2@�q�q�?             @        ������������������������       �                     @                              03C7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 @(;L]n�?             >@                                 �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ;@        	                         @X�<ݚ�?             2@       
                         �?��.k���?             1@                              ���X@և���X�?             @        ������������������������       �                     @                              �̒f@      �?             @                             `f^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                �B@���Q��?             $@                                ,@�q�q�?             @        ������������������������       �                      @                              �̾w@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������Q�Ȟ���?^-n����?X9��v��?���Mb�?|���?|���?      �?        ձ�6Ls�?qBJ�eD�?W�+�ɕ?}g���Q�?UUUUUU�?�������?      �?      �?              �?      �?                      �?              �?�a�a�?��<��<�?UUUUUU�?�������?              �?h/�����?�Kh/��?UUUUUU�?�������?              �?      �?        �a�a�?��y��y�?      �?                      �?              �?�V'u�?��}ylE�?      �?      �?      �?      �?              �?      �?        �$I�$I�?�m۶m��?F]t�E�?]t�E�?              �?�������?�������?      �?      �?      �?      �?              �?      �?                      �?              �?              �?6eMYS��?�5eMYS�?�q�q�?9��8���?              �?�������?333333�?              �?      �?      �?      �?      �?              �?      �?              �?      �?      �?                      �?(�Y�	q�?�wL��?      �?        ------�?�������?              �?�E]t��?]t�E]�?G}g����?r1����?�0�0�?z��y���?��؉���?ى�؉��?      �?        UUUUUU�?�������?]t�E�?F]t�E�?�������?UUUUUU�?�������?�������?      �?              �?      �?      �?                      �?      �?              �?        vb'vb'�?;�;��?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?      �?�$I�$I�?۶m۶m�?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ���@���?Y��"��?ߚ�Cq��?����:.�?�������?�������?�v%jW��?��+Q��?�Y7�"��?L�Ϻ��?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?ى�؉��?�؉�؉�?�������?UUUUUU�?xxxxxx�?�?      �?        UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?              �?                      �?      �?        �������?UUUUUU�?      �?        �؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��\�?���G'�?�Y�"�?�3�뎷?UUUUUU�?UUUUUU�?      �?                      �?����9�?�g�#1�?�̻���?.�!J粹?9��8���?�q�q�?      �?        $�;��?qG�w��?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?      �?                      �?��{a�?a���{�?�z�G��?{�G�z�?�������?UUUUUU�?      �?        �m۶m��?�$I�$I�?      �?        333333�?�������?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        蝺����?�+J�#�?�\AL� �?x6�;��?UUUUUU�?UUUUUU�?      �?        �������?�������?��Moz��?Y�B��?=��<���?�a�a�?      �?              �?      �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?        �5��P�?(�����?���{��?�B!��?      �?              �?      �?              �?      �?        Sa���i�?���!pc�?��[��[�?�A�A�?��4>2��?�Ե��?�V'u�?'u_[�?|���?|���?UUUUUU�?UUUUUU�?      �?              �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?333333�?�������?      �?                      �?8��18�?������?      �?              �?      �?��{���?�B!��?      �?      �?      �?              �?      �?      �?              �?        �������?�������?              �?      �?              �?        ��؉���?ى�؉��?UUUUUU�?�������?�k(���?(�����?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?        �������?333333�?      �?      �?              �?      �?              �?      �?      �?        ?�>��?l�l��?              �?F]t�E�?F]t�E�?�Mozӛ�?d!Y�B�?��8��8�?�q�q�?      �?        �������?�������?      �?      �?      �?              �?      �?      �?              �?              �?              �?      �?      �?      �?UUUUUU�?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�?UUUUUU�?UUUUUU�?              �?      �?              �?        r�q��?�q�q�?�������?�?۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?      �?                      �?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJnխphG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM)hjh))��}�(h,h/h0M)��h2h3h4hph<�h=Kub������       \                    �?<C�`��?�           8�@               S                    @��1+�?�            �m@              R                    @F����?�            �k@              E                   �E@(w's�M�?�            �j@                                   @r ��*�?t            �g@                                  �?`'�J�?@            �Y@        ������������������������       �                     ;@                                   �?Х-��ٹ?.            �R@       	                          @0@�i�y�?&            �O@        
                          �B@؇���X�?	             ,@                                 �9@$�q-�?             *@                                  �6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                    �H@                                   @r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@                                 ��@�^�����?4            �U@                                �|Y:@�+$�jP�?             ;@                               ��@�IєX�?             1@       ������������������������       �                     (@                                  �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                �&�@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @               ,                    �?:���W�?'            �M@                !                    3@ �o_��?             9@        ������������������������       �                     $@        "       #                    �?��S���?	             .@        ������������������������       �                     @        $       %                   �7@�z�G��?             $@        ������������������������       �                     @        &       +                    �?      �?             @       '       *                  SE"@���Q��?             @       (       )                 �|Y>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        -       8                    �?j���� �?             A@        .       7                    �?�<ݚ�?             2@       /       6                  S�-@�	j*D�?             *@        0       5                 ���,@�q�q�?             @       1       2                 �&�)@�q�q�?             @        ������������������������       �                     �?        3       4                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        9       :                 P��%@      �?             0@        ������������������������       �                     @        ;       D                    �?      �?
             (@       <       =                    &@���Q��?             $@        ������������������������       �                     @        >       ?                 �|�7@և���X�?             @        ������������������������       �                     @        @       A                    �?      �?             @        ������������������������       �                      @        B       C                   �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        F       Q                 `f~B@R�}e�.�?             :@        G       L                    �?�q�q�?             (@       H       I                    (@�q�q�?             @        ������������������������       �                     �?        J       K                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        M       P                   P>@r�q��?             @       N       O                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        ������������������������       �                     "@        T       U                   -@      �?             0@        ������������������������       �                     �?        V       W                    �?��S�ۿ?             .@        ������������������������       �                     @        X       [                    @�8��8��?	             (@        Y       Z                 ff.b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ]                       Ј�U@�:�B��?(           �}@       ^       �                    �?��S�sT�?           P|@        _       �                    �?p�}�ޤ�?0            @R@       `       o                     @L=�m��?'            �N@        a       b                 ���=@؇���X�?             5@        ������������������������       �                     @        c       n                   �M@d}h���?	             ,@       d       k                    �?�z�G��?             $@       e       j                 `f�A@      �?              @       f       g                  Y>@�q�q�?             @        ������������������������       �                     �?        h       i                 X�lA@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        l       m                     �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        p                           �?z�G�z�?             D@       q       ~                 @3s+@�<ݚ�?             B@       r       s                   �6@@�0�!��?             A@        ������������������������       �                     @        t       u                 ���@��a�n`�?             ?@        ������������������������       �                     &@        v       }                 �|�=@R���Q�?             4@       w       x                   �<@z�G�z�?             .@        ������������������������       �                     @        y       z                   @@      �?             (@        ������������������������       �      �?              @        {       |                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?	             (@        �       �                    F@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 ��y&@���Q��?             @        ������������������������       �                     �?        �       �                     @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��$:@X�����?�            �w@       �       �                  ��@����-��?�            �q@        ������������������������       �        %             O@        �       �                    �?���,��?�            �k@       �       �                    �?�7��t�?�            �j@        �       �                   `3@؇���X�?             <@       �       �                 �|Y=@�����H�?             ;@        ������������������������       �                      @        �       �                    �?`2U0*��?             9@       �       �                 ��(@      �?
             0@       �       �                 X��A@�C��2(�?             &@       ������������������������       ������H�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?0�#�.^�?            `g@       �       �                     @�(̶h�?z            @f@        �       �                    �?��S�ۿ?&             N@       �       �                    4@����˵�?%            �M@        �       �                   �2@"pc�
�?             &@        ������������������������       �                     @        �       �                   �'@����X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        �       �                     �?@��8��?             H@        ������������������������       �                     @        �       �                    �?`���i��?             F@       �       �                   �@@�?�|�?            �B@        ������������������������       �                     5@        �       �                   @A@      �?             0@        ������������������������       ��q�q�?             @        ������������������������       �        	             *@        ������������������������       �                     @        ������������������������       �                     �?        �       �                    )@��g�g�?T            �]@        ������������������������       �                      @        �       �                 ��) @��Õty�?S             ]@       �       �                    �?l{��b��?5            �S@       �       �                 �Yu@$�q-�?4            �S@        �       �                 ��@؇���X�?             5@        ������������������������       �                     @        �       �                 �|�;@@�0�!��?             1@       ������������������������       �                     "@        �       �                 �&B@      �?              @       �       �                 �|Y>@����X�?             @        ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �>@�}�+r��?&            �L@       �       �                 @3�@p���?             I@        ������������������������       �                     8@        �       �                   �1@ ��WV�?             :@        ������������������������       �r�q��?             @        ������������������������       �                     4@        �       �                   �?@����X�?             @        ������������������������       �                     �?        �       �                   @C@r�q��?             @       ������������������������       �                     @        �       �                   �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    9@��G���?            �B@        ������������������������       �                     "@        �       �                    �?      �?             <@       �       �                   �;@�q�q�?             8@        ������������������������       �                      @        �       �                    �?�GN�z�?             6@       �       �                   �<@�d�����?             3@        ������������������������       �                     @        �       �                   @A@X�Cc�?
             ,@       �       �                    (@�eP*L��?             &@       �       �                 `��!@      �?              @        ������������������������       �                      @        �       �                 �|�=@      �?             @       �       �                 ���"@      �?             @        ������������������������       �                      @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                 ��I7@����X�?             @       �       �                    +@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �                          R@      �?7             X@       �                          �?��<b���?6             W@       �                          �?�1�`jg�?             �K@       �       �                   �>@l��
I��?             K@       �       �                    D@l��[B��?             =@        �       �                   �<@d}h���?             ,@        ������������������������       �                     @        �       �                 03k:@�z�G��?             $@        ������������������������       �                     @        �       �                   @>@և���X�?             @       �       �                 `fF<@���Q��?             @        �       �                 �|�?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �J@z�G�z�?             .@        �       �                    H@      �?              @       �       �                   �F@r�q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �                          ;@HP�s��?             9@                                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   @�nkK�?             7@       ������������������������       �                     5@                              �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        	                         @������?            �B@        
                         @      �?             @                                @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                 �?�FVQ&�?            �@@        ������������������������       �                      @                                  �?`Jj��?             ?@                              ��9L@�t����?             1@       ������������������������       �                     &@                              03�M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             ,@        ������������������������       �                     @              $                ���a@p�ݯ��?
             3@             #                   �?"pc�
�?             &@                                �?�<ݚ�?             "@                                �B@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?              "                   �?      �?             @              !                @�pX@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        %      (                   �?      �?              @       &      '                �̾w@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0M)KK��h2h3h4hVh<�h=Kub�������������܍�W�?/�F�JP�?0]�X#�?hQ�Sn��?;Ӹ�Qg�?1ˑ�+f�?]���~!�?)��L�w�?R�٨�l�?,�����?�?�������?              �?O贁N�?K~��K�?AA�?�������?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?      �?                      �?UUUUUU�?�������?      �?                      �?֔5eMY�?�5eMYS�?B{	�%��?/�����?�?�?              �?�������?�������?      �?                      �?�������?333333�?      �?                      �?A�Iݗ��?_[4��?�Q����?
ףp=
�?              �?�������?�?              �?ffffff�?333333�?      �?              �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?ZZZZZZ�?�������?�q�q�?9��8���?;�;��?vb'vb'�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?              �?      �?      �?      �?              �?      �?�������?333333�?              �?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        �;�;�?'vb'vb�?�������?�������?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?              �?      �?              �?�������?�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �c+����?�pR���?/��K2�?D�L�6�?�z��ի�?�
*T��?���:�?�����?۶m۶m�?�$I�$I�?      �?        I�$I�$�?۶m۶m�?ffffff�?333333�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?      �?              �?      �?              �?        �������?�������?9��8���?�q�q�?ZZZZZZ�?�������?              �?�s�9��?�c�1Ƹ?      �?        333333�?333333�?�������?�������?      �?              �?      �?      �?      �?      �?      �?              �?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?�$I�$I�?�m۶m��?              �?      �?        �������?333333�?      �?              �?      �?      �?                      �?�=�ĩ��?#�X��?ܥ���.�? �
���?      �?        X��;ze�?C�I .Լ?X:Ɂ���??-���b�?۶m۶m�?�$I�$I�?�q�q�?�q�q�?              �?���Q��?{�G�z�?      �?      �?]t�E�?F]t�E�?�q�q�?�q�q�?      �?              �?              �?                      �?��b���?w��?�JV����?��MmjS�?�������?�?W'u_�?��/���?/�袋.�?F]t�E�?      �?        �m۶m��?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?        F]t�E�?F]t�E�?*�Y7�"�?к����?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?                      �?ي����?��}ylE�?              �?�FX�i�?��=���?${�ґ�?�&��jq�?�؉�؉�?;�;��?۶m۶m�?�$I�$I�?      �?        ZZZZZZ�?�������?      �?              �?      �?�m۶m��?�$I�$I�?333333�?�������?      �?                      �?�5��P�?(�����?\���(\�?{�G�z�?      �?        O��N���?;�;��?�������?UUUUUU�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?        #�u�)��?v�)�Y7�?      �?              �?      �?�������?�������?              �?�袋.��?]t�E�?Cy�5��?y�5���?      �?        %I�$I��?�m۶m��?t�E]t�?]t�E�?      �?      �?              �?      �?      �?      �?      �?      �?              �?      �?              �?      �?                      �?      �?              �?              �?              �?              �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?��,d!�?��Moz��?��k߰�?��)A��?Lh/����?h/�����?���=��?GX�i���?۶m۶m�?I�$I�$�?              �?333333�?ffffff�?              �?۶m۶m�?�$I�$I�?333333�?�������?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        q=
ףp�?{�G�z�?      �?      �?      �?                      �?�Mozӛ�?d!Y�B�?      �?              �?      �?      �?                      �?      �?        ��g�`��?к����?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?>����?|���?      �?        ���{��?�B!��?<<<<<<�?�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?Cy�5��?^Cy�5�?F]t�E�?/�袋.�?�q�q�?9��8���?�������?�������?              �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?�$I�$I�?۶m۶m�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�[�.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       b                    �?�,�٧��?�           8�@                                `f�%@0�".���?�            �p@                                �̌@      �?"             J@                                   �?"pc�
�?             6@                               �|�9@      �?             0@        ������������������������       �                     @                                ���@z�G�z�?             $@        ������������������������       �                     �?        	       
                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?                                ���@�q�q�?             @        ������������������������       �                     �?                                   4@���Q��?             @        ������������������������       �                     �?                                pf�@      �?             @                               �|Y:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                    @������?             >@                                  �J@      �?              @       ������������������������       �                     @        ������������������������       �                      @                                   3@�C��2(�?             6@        ������������������������       �                     �?                                �|Y>@���N8�?
             5@       ������������������������       �        	             4@        ������������������������       �                     �?               G                    �?]���?�             k@              @                 Ь�9@�5U��K�?h            �d@                %                    �?     ��?1             T@        !       "                 P�>,@�?�|�?            �B@       ������������������������       �                     =@        #       $                 pF4.@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        &       ?                   �D@��V#�?            �E@       '       >                  ��8@��i#[�?             E@       (       ;                 `v�5@������?            �D@       )       0                 �|�<@     ��?             @@       *       /                    @��.k���?             1@       +       ,                 �B,@X�Cc�?
             ,@        ������������������������       �                     @        -       .                   �0@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        1       :                    @@z�G�z�?
             .@       2       3                  S�-@      �?             (@        ������������������������       �                      @        4       5                    �?ףp=
�?             $@        ������������������������       �                     @        6       7                 ��1@r�q��?             @        ������������������������       �                     @        8       9                 03C3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        <       =                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        A       F                    :@��f�{��?7            �U@        B       C                    �?�C��2(�?             &@        ������������������������       �                     @        D       E                   �E@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        /            �R@        H       Q                    �?j���� �?"            �I@        I       P                    �?�����?             5@        J       O                  18@      �?              @       K       N                    @؇���X�?             @       L       M                 �|Y=@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        R       S                    �?d��0u��?             >@        ������������������������       �                     @        T       W                    @l��
I��?             ;@        U       V                    @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        X       Y                 ��5@�GN�z�?             6@        ������������������������       �                     �?        Z       [                     @��s����?             5@        ������������������������       �                     @        \       ]                    @�X�<ݺ?             2@       ������������������������       �        
             .@        ^       _                 ��T?@�q�q�?             @        ������������������������       �                     �?        `       a                 pf�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        c       �                 ��%@�
8\��?           �{@       d       u                    �?l�b�G��?�            �l@        e       r                    �?PN��T'�?             ;@       f       g                   �7@�LQ�1	�?             7@        ������������������������       �                     �?        h       k                 �|Y=@�C��2(�?             6@        i       j                   @@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        l       q                 X�,@@�IєX�?	             1@       m       p                   @@@4և���?             ,@       n       o                 ���@ףp=
�?             $@        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        s       t                 ��}@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        v       w                 ���@�L#���?�             i@        ������������������������       �                     9@        x       �                    �?t��ճC�?q             f@       y       ~                    �?l�b�G��?n            `e@        z       }                 �|Y=@�KM�]�?
             3@        {       |                  ��@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     .@               �                   �3@`-�I�w�?d             c@        �       �                 �?�@���y4F�?             3@        ������������������������       �                     $@        �       �                 pf� @X�<ݚ�?             "@        �       �                   �1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 ���@P#aE�?V            �`@        ������������������������       �                      @        �       �                   �:@ ����O�?U            ``@        ������������������������       �                     E@        �       �                     @ p�/��?8            @V@        ������������������������       �                     @        �       �                 @Q!@��`qM|�?4            �T@       �       �                 @3�@      �?,             P@       �       �                   �?@���N8�?             E@       ������������������������       �                     9@        �       �                   �E@�t����?
             1@       �       �                   �B@z�G�z�?             $@       �       �                 �&B@�����H�?             "@        ������������������������       �                     @        �       �                 P�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     6@        �       �                   �;@�KM�]�?             3@        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     @        �                        @�:x@�X�2�?�            �j@       �       �                 �&@�s5��&�?�            @j@        ������������������������       �                      @        �       �                    @~e�.y��?�             j@        �       �                     @��Q��?             4@        ������������������������       �                     $@        �       �                    �?�z�G��?             $@        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     @        �       �                 ��T?@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @ظ�*���?y            �g@       �       �                     �?6�h_�?u            �f@        �       �                 �\@<�\`*��?3             U@       �       �                    �?:%�[��?,            �Q@       �       �                    �?=��T�?+            �Q@       �       �                   �J@θ	j*�?             J@       �       �                  �>@��.k���?             A@        �       �                 �|�?@�t����?
             1@       �       �                   @>@�eP*L��?             &@       �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                 `f�;@r�q��?             @        ������������������������       �                      @        �       �                 �|Y=@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 `��L@������?             1@       �       �                   �B@     ��?             0@        �       �                 X�lA@�q�q�?             "@       �       �                 �|�<@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�X�<ݺ?	             2@       �       �                    �?@4և���?             ,@        ������������������������       �                     @        �       �                   �Q@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?X�<ݚ�?             2@        ������������������������       �                     @        �       �                  x#J@�q�q�?             (@        ������������������������       �                      @        �       �                    �?���Q��?             $@       �       �                 `�iJ@X�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?����X�?             @       �       �                 03�Q@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?$�q-�?             *@        �       �                 X��C@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    $@�C��2(�?B            �X@        ������������������������       �                      @        �       �                   �A@,���$�?A            @X@       �       �                   �@@H�ՠ&��?)             K@       �       �                    �?4��?�?(             J@        �       �                    �?d}h���?             ,@       �       �                     @ףp=
�?	             $@        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �y_:@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �9@�}�+r��?             C@       ������������������������       �                     2@        �       �                   �:@ףp=
�?             4@        �       �                  �DC@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�=@�X�<ݺ?             2@       �       �                   �+@�8��8��?             (@        �       �                 �|Y<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �E@        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������&��jq�?:�g *�?�� ;J��?�?qm��?      �?      �?F]t�E�?/�袋.�?      �?      �?              �?�������?�������?      �?        �q�q�?�q�q�?              �?      �?        UUUUUU�?UUUUUU�?              �?�������?333333�?      �?              �?      �?      �?      �?              �?      �?                      �?wwwwww�?�?      �?      �?              �?      �?        ]t�E�?F]t�E�?              �?��y��y�?�a�a�?      �?                      �?�LW�+��?�,j5��?��k���?���h��?      �?      �?к����?*�Y7�"�?              �?      �?      �?      �?                      �?6eMYS��?eMYS֔�?�<��<��?�a�a�?��+Q��?�v%jW��?      �?      �?�?�������?�m۶m��?%I�$I��?              �?]t�E�?t�E]t�?              �?      �?              �?        �������?�������?      �?      �?      �?        �������?�������?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?�q�q�?              �?      �?              �?              �?        �}A_Ї?������?F]t�E�?]t�E�?              �?�$I�$I�?۶m۶m�?              �?      �?                      �?ZZZZZZ�?�������?�a�a�?=��<���?      �?      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?                      �?DDDDDD�?wwwwww�?              �?Lh/����?h/�����?�������?333333�?      �?                      �?�袋.��?]t�E�?              �?z��y���?�a�a�?              �?��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �����?��#��#�?�Gp��?p�}��?&���^B�?h/�����?��Moz��?Y�B��?              �?]t�E�?F]t�E�?�������?�������?      �?                      �?�?�?n۶m۶�?�$I�$I�?�������?�������?      �?              �?      �?      �?              �?              �?      �?      �?                      �?��@���?g��1��?      �?        �E]t��?t�E]t�?�Gp��?p�}��?�k(���?(�����?      �?      �?      �?                      �?      �?        Q^Cy��?y�5�װ?6��P^C�?(������?      �?        r�q��?�q�q�?      �?      �?      �?                      �?�������?�������?      �?      �?      �?        �蛣o��?�qA��?              �?����?qBJ�eD�?      �?        �G?�я�?p�\��?      �?        �@	o4u�?��k���?      �?      �?��y��y�?�a�a�?      �?        <<<<<<�?�?�������?�������?�q�q�?�q�q�?      �?        �������?�������?              �?      �?                      �?      �?              �?        �k(���?(�����?              �?      �?              �?        ����z�?�Zn��?�~��~��?p'p'�?              �?vb'vb'�?'vb'vb�?ffffff�?�������?              �?ffffff�?333333�?      �?              �?      �?      �?        �������?333333�?      �?                      �?&W�+��?g���Q��?��o��Z�?�Y@�H��?=��<���?�a�a�?+l$Za�?�'�K=�?�:��:��?�������?�؉�؉�?�N��N��?�������?�?�������?�������?]t�E�?t�E]t�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?      �?                      �?              �?              �?xxxxxx�?�?      �?      �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?                      �?      �?                      �?��8��8�?�q�q�?n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?      �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?        333333�?�������?r�q��?�q�q�?              �?�m۶m��?�$I�$I�?333333�?�������?      �?                      �?      �?              �?                      �?�؉�؉�?;�;��?�������?�������?      �?                      �?      �?        ]t�E�?F]t�E�?              �?�,O"Ӱ�?���fy�?������?{	�%���?�N��N��?ى�؉��?I�$I�$�?۶m۶m�?�������?�������?      �?        �������?UUUUUU�?      �?                      �?      �?      �?              �?      �?        �5��P�?(�����?      �?        �������?�������?      �?      �?      �?                      �?��8��8�?�q�q�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?      �?              �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��=hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM7hjh))��}�(h,h/h0M7��h2h3h4hph<�h=Kub������       |                     @���*1�?�           8�@               W                   @K@���0��?�            @t@              &                    �?\I�~�?�            �l@               	                    �?H0sE�d�?/            �R@                                    �?8�Z$���?             *@                                  �H@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        
       %                    :@��a�n`�?)             O@              $                   �J@"pc�
�?            �@@              #                    G@     ��?             @@              "                   �E@�q�q�?             8@                                 �6@��2(&�?             6@        ������������������������       �                     @                                  �;@z�G�z�?             .@                                  �9@      �?             @                                  �?�q�q�?             @                                 �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?               !                    �?�C��2(�?	             &@                                  �?      �?              @        ������������������������       �                     �?                                  �'@؇���X�?             @        ������������������������       �                     �?                                  �A@r�q��?             @       ������������������������       �                     @                                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     =@        '       (                    #@Tݭg_�?]            �c@        ������������������������       �                     $@        )       F                     �?��ӄ���?X            @b@        *       A                    �?      �?'             N@       +       @                    �?R�}e�.�?#             J@       ,       -                   �<@t�F�}�?"            �I@        ������������������������       �                     @        .       ?                   �>@�3Ea�$�?             G@       /       0                 `fF:@8�A�0��?             6@        ������������������������       �                     @        1       <                 ���=@      �?             2@       2       ;                   @K@և���X�?             ,@       3       :                    @@���Q��?             $@        4       9                    �?z�G�z�?             @       5       8                 �|�=@�q�q�?             @       6       7                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        =       >                   @D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     8@        ������������������������       �                     �?        B       E                 `�iJ@      �?              @        C       D                  x#J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        G       V                   �*@ �#�Ѵ�?1            �U@       H       I                    �?�NW���?            �J@        ������������������������       �                      @        J       K                    @�:�]��?            �I@        ������������������������       �                      @        L       U                 �|�=@�ʈD��?            �E@       M       T                    �?"pc�
�?             6@       N       S                 �|�<@�<ݚ�?             2@       O       R                    5@      �?
             0@        P       Q                    &@����X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@        ������������������������       �                    �@@        X       m                   �E@r֛w���?;            @W@       Y       ^                    �?�~t��?/            @Q@       Z       [                    �?�&=�w��?#            �J@       ������������������������       �                     F@        \       ]                    $@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        _       h                 �|Y>@      �?             0@       `       g                    �?���|���?             &@       a       b                   �7@      �?              @        ������������������������       �                      @        c       f                    �?�q�q�?             @        d       e                 0c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        i       l                    �?z�G�z�?             @        j       k                 pU�t@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        n       u                   �I@�q�q�?             8@        o       p                   �G@"pc�
�?             &@        ������������������������       �                     @        q       t                    �?�q�q�?             @        r       s                 �UkT@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        v       w                    �?�n_Y�K�?             *@        ������������������������       �                     @        x       y                    �?�����H�?             "@        ������������������������       �                     @        z       {                   �T@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        }       �                 P��%@���t�?�            0x@       ~       �                 �̌@^wUBO��?�            �m@              �                    �?�i��D�?N            �`@        �       �                 `�j@F�����?&            @R@       �       �                   �6@�t����?$             Q@        �       �                    �?�z�G��?             $@       �       �                    �?�<ݚ�?             "@       �       �                    �?      �?              @        ������������������������       �                     �?        �       �                 ��y@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?^l��[B�?             M@       �       �                    �?�MWl��?            �L@        �       �                 ���@      �?             (@        ������������������������       �                     �?        �       �                  s�@"pc�
�?             &@        ������������������������       �                      @        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                 ���@�:�^���?            �F@        ������������������������       �                     (@        �       �                 ���@<���D�?            �@@        �       �                 �|�:@����X�?             @        ������������������������       �                     �?        �       �                 �|�=@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        �       �                 ���@$�q-�?             :@        ������������������������       �                     @        �       �                 ��(@�KM�]�?	             3@       �       �                 X�I@�����H�?             2@       ������������������������       ��r����?             .@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���*�?(             N@       �       �                    ;@F�4�Dj�?'            �M@       �       �                    �?      �?             @@        �       �                 �&B@      �?              @       �       �                 ���@      �?             @        ������������������������       �                      @        �       �                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �? �q�q�?             8@       �       �                    7@�nkK�?             7@       ������������������������       �        
             ,@        �       �                   �8@�����H�?             "@        �       �                 �&b@      �?             @        ������������������������       �                      @        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 pf�@�����H�?             ;@       ������������������������       �        
             1@        �       �                   �?@�z�G��?             $@       �       �                 �|Y=@      �?              @        ������������������������       �                     @        �       �                 �|Y>@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �?�@���C��?J            �Z@        ������������������������       �                     7@        �       �                   @9@���O1��?7            �T@        �       �                   �2@��p\�?            �D@        �       �                 @�"@8�Z$���?             *@       �       �                 ��Y @�8��8��?             (@        �       �                    1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?h�����?             <@        ������������������������       �                     @        �       �                    �?���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        �       �                 ��) @d}h���?             E@       �       �                 @3�@ �Cc}�?             <@        �       �                   �?@���Q��?             @        ������������������������       �                      @        �       �                   �A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        �       �                    �?և���X�?	             ,@        ������������������������       �                     �?        �       �                    �?��
ц��?             *@       �       �                 �|�>@      �?             (@       �       �                   `!@�q�q�?             "@        ������������������������       �                     @        �       �                   �<@���Q��?             @        ������������������������       �                      @        �       �                 `f6"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �                       03�7@rr�J��?X            �b@       �                         �?@���L��?6            �V@       �                          �?��c�%�?/            @S@       �       �                 ��*@�j�'�=�?(            �P@        ������������������������       �                     &@        �       �                    @�b��[��?"            �K@        ������������������������       �                     @        �       �                 `�X.@Fx$(�?              I@        �       �                    �?�<ݚ�?             "@        �       �                    �?���Q��?             @       �       �                   �-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �                          �?������?            �D@       �                           �?�>4և��?             <@       �       �                   �0@R���Q�?             4@        ������������������������       �                     �?        �       �                 ��.@�KM�]�?             3@        �       �                 �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     .@                                 �?      �?              @                              �|�;@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                �0@��
ц��?             *@        ������������������������       �                      @                                 �?���|���?
             &@       	                         �?և���X�?             @       
                      ��1@���Q��?             @                             �|�;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                               �v6@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @                                @C@@4և���?             ,@                                 �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @              "                   �?���5��?"            �L@              !                   �?և���X�?             @                             �T)D@      �?             @        ������������������������       �                      @                                 ;@      �?             @        ������������������������       �                      @                                  >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        #      6                   @HP�s��?             I@       $      %                   �?�����?             E@        ������������������������       �                     @        &      '                   �?�KM�]�?             C@        ������������������������       �                     (@        (      1                   @8�Z$���?             :@       )      *                   @z�G�z�?	             .@        ������������������������       �                     @        +      0                   �?�q�q�?             "@       ,      /                   @      �?              @        -      .                   @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        2      3                ��T?@�C��2(�?             &@        ������������������������       �                      @        4      5                ���A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0M7KK��h2h3h4hVh<�h=Kub������������`l����??'��d�?���Kh�?����K�?!��O���?�cj`��?O贁N�?��b�/��?;�;��?;�;��?      �?      �?              �?      �?                      �?�c�1Ƹ?�s�9��?F]t�E�?/�袋.�?      �?      �?�������?UUUUUU�?t�E]t�?��.���?              �?�������?�������?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?        F]t�E�?]t�E�?      �?      �?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?      �?                      �?� � �?�|˷|��?              �?_�z����?�
*T��?      �?      �?'vb'vb�?�;�;�?777777�?�������?              �?����7��?��,d!�?颋.���?/�袋.�?      �?              �?      �?�$I�$I�?۶m۶m�?�������?333333�?�������?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?      �?              �?      �?      �?                      �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �/����?�}A_Ч?萚`���?�x+�R�?      �?        }}}}}}�?�?      �?        A_���?�}A_з?/�袋.�?F]t�E�?9��8���?�q�q�?      �?      �?�m۶m��?�$I�$I�?      �?      �?      �?              �?                      �?      �?              �?              �?        �B!��?���{��?)�3J���?�s��\�?�x+�R�?tHM0���?              �?�q�q�?9��8���?      �?                      �?      �?      �?]t�E]�?F]t�E�?      �?      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        ى�؉��?;�;��?      �?        �q�q�?�q�q�?              �?      �?      �?      �?                      �?�mF2<�?b$�s���?�=����?M�[��?ju�՝V�?,�T�R�?�P�B�
�?�^�z���?�������?�������?333333�?ffffff�?�q�q�?9��8���?      �?      �?              �?�$I�$I�?�m۶m��?      �?                      �?              �?      �?        �=�����?��=���?:��,���?�YLg1�?      �?      �?      �?        F]t�E�?/�袋.�?              �?�q�q�?9��8���?              �?      �?        }�'}�'�?l�l��?      �?        |���?|���?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?        �؉�؉�?;�;��?      �?        �k(���?(�����?�q�q�?�q�q�?�������?�?      �?              �?              �?                      �?""""""�?wwwwww�?��/���?�A�I��?      �?      �?      �?      �?      �?      �?              �?      �?      �?      �?                      �?              �?�������?UUUUUU�?�Mozӛ�?d!Y�B�?      �?        �q�q�?�q�q�?      �?      �?      �?              �?      �?              �?      �?              �?              �?        �q�q�?�q�q�?      �?        ffffff�?333333�?      �?      �?      �?        �������?�������?      �?      �?      �?                      �?      �?        \�琚`�?"5�x+��?      �?        P�M�_�?���ˊ��?�]�ڕ��?��+Q��?;�;��?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�m۶m��?�$I�$I�?      �?        �.�袋�?F]t�E�?      �?                      �?I�$I�$�?۶m۶m�?%I�$I��?۶m۶m�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?        �;�;�?�؉�؉�?      �?      �?UUUUUU�?UUUUUU�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        Z7�"�u�?L�Ϻ��?�!�!�?�����?(�Y�	q�?�S{��?m��&�l�?�&�l���?              �?־a��?� O	��?              �?R���Q�?ףp=
��?9��8���?�q�q�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ��+Q��?�v%jW��?�m۶m��?�$I�$I�?333333�?333333�?      �?        (�����?�k(���?      �?      �?              �?      �?                      �?      �?      �?�������?333333�?              �?      �?                      �?�;�;�?�؉�؉�?              �?]t�E]�?F]t�E�?۶m۶m�?�$I�$I�?333333�?�������?      �?      �?      �?                      �?      �?                      �?      �?        F]t�E�?t�E]t�?      �?                      �?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?              �?      �?              �?        �}��?��Gp�?�$I�$I�?۶m۶m�?      �?      �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        q=
ףp�?{�G�z�?=��<���?�a�a�?      �?        �k(���?(�����?      �?        ;�;��?;�;��?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?                      �?      �?                      �?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��(hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                    �?n��"�)�?�           8�@              A                    �?(��g���?a           8�@                                    �?P�;�&��?d            @e@                                   �?�nkK�?%            @Q@                                 �H@�L���?            �B@       ������������������������       �                     ?@               
                    �?      �?             @              	                    K@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @@               @                    �?N��>��??            @Y@                                   @      �?>             Y@                                  �&@��G���?            �B@                                  �J@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @                                  �,@      �?             @@                                   �?������?
             1@        ������������������������       �                      @                                  �B@������?             .@                               `f�)@�C��2(�?             &@        ������������������������       �                      @                                   ;@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                                   D@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             .@                )                    �?����X�?'            �O@        !       (                    �? ��WV�?             :@        "       #                    �?      �?             @        ������������������������       �                     �?        $       %                 �&�)@�q�q�?             @        ������������������������       �                     �?        &       '                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        *       ?                   @B@��%��?            �B@       +       6                   �6@      �?             @@        ,       1                 xF� @�q�q�?	             (@        -       .                 ���@      �?             @        ������������������������       �                     �?        /       0                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        2       5                    �?      �?              @       3       4                  �#@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        7       >                 ��� @z�G�z�?
             4@       8       =                    ;@���|���?             &@       9       <                   �9@      �?              @        :       ;                 pf�@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     �?        B       �                 ���=@ĩ����?�            �w@       C       �                   @E@XT�z�q�?�            �s@       D       I                     �?�p�Ð�?�            Pq@        E       F                    �?����X�?             ,@        ������������������������       �                      @        G       H                 �|�<@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        J       �                   @C@�ɱK���?�            pp@       K       L                 ���@��k�c��?�            `o@        ������������������������       �                     8@        M       N                 ��@�E���?�            `l@        ������������������������       �                      @        O       T                  ��@H0sE�d�?�             l@        P       S                 �Y�@ ��WV�?             :@        Q       R                 ���@ףp=
�?             $@       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     0@        U       Z                 ��@P���+�?�            �h@        V       W                 �|Y=@���!pc�?             &@        ������������������������       �                     �?        X       Y                    �?z�G�z�?             $@       ������������������������       �      �?              @        ������������������������       �                      @        [       j                   �4@�*/�8V�?|            �g@        \       c                 ��Y @:�&���?            �C@        ]       ^                 �?�@      �?             0@       ������������������������       �                      @        _       `                 @3�@      �?              @        ������������������������       �                      @        a       b                   �1@�q�q�?             @        ������������������������       �      �?              @        ������������������������       �      �?             @        d       e                 `�X$@�nkK�?             7@        ������������������������       �                     (@        f       g                   �2@�C��2(�?             &@       ������������������������       �                      @        h       i                   �'@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        k       �                    �?�
�@c�?a            �b@       l       �                   �>@R�xE��?Q            �_@       m       t                     @���1j	�?:            �U@        n       o                 �|�<@      �?             0@       ������������������������       �                     $@        p       s                 �|�=@r�q��?             @        q       r                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        u       �                 �|Y=@ >�֕�?/            �Q@        v                          �<@�t����?             A@       w       x                    �?     ��?             @@        ������������������������       �                      @        y       z                 pf� @(;L]n�?             >@       ������������������������       �                     4@        {       ~                 @3"@ףp=
�?             $@        |       }                    8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     B@        �       �                    �?��r._�?            �D@        ������������������������       �                     @        �       �                   �?@>A�F<�?             C@        �       �                 pff@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     @؇���X�?            �A@        �       �                   �@@      �?              @        ������������������������       �                      @        �       �                   �A@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        �       �                   �@�����H�?             ;@        �       �                   @@@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @@@�nkK�?             7@        �       �                 ��I @�����H�?             "@       ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     ,@        �       �                    �?���7�?             6@        �       �                  �v6@�����H�?             "@       ������������������������       �                     @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             *@        �       �                    �?�q�q�?	             (@       �       �                   �C@X�<ݚ�?             "@        �       �                     @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     @�q�q�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �D@        �       �                    �?�G��l��?*            �O@       �       �                 �!fK@П[;U��?(             M@       �       �                    �?ҳ�wY;�?             A@       �       �                    �?�f7�z�?             =@        �       �                 �|�;@և���X�?             @        ������������������������       �                      @        �       �                 X�lA@z�G�z�?             @        ������������������������       �                      @        �       �                 p�i@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �<@8�A�0��?             6@        �       �                 `f�D@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �H@�q�q�?             2@       �       �                 X�,C@r�q��?             (@       �       �                   �>@�<ݚ�?             "@        �       �                 �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 03�D@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 p"�X@�q�q�?             8@       �       �                   �8@������?             1@        ������������������������       �                     �?        �       �                      @     ��?             0@       �       �                   �D@�8��8��?             (@       ������������������������       �                     @        �       �                 ЈT@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    ;@      �?             @        ������������������������       �                     �?        �       �                 �|�>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 p�w@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �                          @H�z�G�?b             d@       �       �                    �?�e����?^            �c@       �       �                    �?4�{Y���?3            �T@       �       �                     @HP�s��?             I@       ������������������������       �                    �@@        �       �                    @������?             1@       �       �                    �?�r����?	             .@        �       �                 �|�7@      �?             @       �       �                   �"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 P��%@�C��2(�?             &@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        �       �                     @:ɨ��?            �@@       ������������������������       �                     3@        �       �                 `f�8@����X�?
             ,@        ������������������������       �                      @        �       �                    @r�q��?	             (@        �       �                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �                          �?X~�pX��?+            @R@       �       �                    )@� �	��?             I@        ������������������������       �        	             ,@        �                            @�<ݚ�?             B@       �       �                    8@؇���X�?             5@        ������������������������       �                      @        �       �                    �?�}�+r��?             3@       �       �                   @B@ףp=
�?             $@        �       �                 @��v@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@                                 �?�q�q�?	             .@                                3@�n_Y�K�?             *@        ������������������������       �                     @                                 �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                 @�nkK�?             7@        	      
                   �?�q�q�?             @        ������������������������       �                     �?                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             4@        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������o怖�?�� 3���?4�[�J	�?��Hej��?�?�������?d!Y�B�?�Mozӛ�?L�Ϻ��?}���g�?              �?      �?      �?333333�?�������?      �?                      �?              �?              �?�tj��?�be�F�?      �?      �?v�)�Y7�?#�u�)��?333333�?�������?              �?      �?              �?      �?�?xxxxxx�?              �?�?wwwwww�?F]t�E�?]t�E�?              �?�q�q�?�q�q�?      �?                      �?      �?      �?      �?                      �?              �?�$I�$I�?�m۶m��?;�;��?O��N���?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?}���g�?���L�?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�������?�������?      �?                      �?      �?        �������?�������?F]t�E�?]t�E]�?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?      �?                      �?�����?`XV��?���3 ��?��c�^�?�U�{�?�gPE!l�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?              �?      �?        ��$�Y�?
��ߖ3�?oI�!m��?���򖄺?      �?        ��z��U�?`�(tSR�?              �?��b�/��?O贁N�?O��N���?;�;��?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?        ���/M�?�Q7���?F]t�E�?t�E]t�?              �?�������?�������?      �?      �?      �?        r1����?m�w6�;�?�A�A�?�o��o��?      �?      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?�Mozӛ�?d!Y�B�?      �?        ]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        �ַC5�?�IA��U�?>������?��`0�?�;⎸#�?qG�wĭ?      �?      �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��+��+�?�A�A�?<<<<<<�?�?      �?      �?              �?�������?�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?              �?        �ڕ�]��?ە�]���?      �?        ������?Cy�5��?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        �q�q�?�q�q�?      �?      �?              �?      �?        �Mozӛ�?d!Y�B�?�q�q�?�q�q�?�������?�������?      �?              �?        �.�袋�?F]t�E�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?r�q��?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?              �?        1�0��?��y��y�?�{a���?��=���?�������?�������?O#,�4��?a���{�?�$I�$I�?۶m۶m�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        颋.���?/�袋.�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?�������?UUUUUU�?9��8���?�q�q�?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?�?xxxxxx�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?�������?�������?      �?                      �?333333�?ffffff�?�A�A�?�-��-��?4u~�!��?�b��7��?{�G�z�?q=
ףp�?              �?�?xxxxxx�?�?�������?      �?      �?      �?      �?              �?      �?                      �?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?      �?        e�M6�d�?N6�d�M�?              �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        �^�z���?�B�
*�?�Q����?)\���(�?              �?9��8���?�q�q�?۶m۶m�?�$I�$I�?              �?�5��P�?(�����?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?;�;��?ى�؉��?      �?        �$I�$I�?�m۶m��?              �?      �?              �?        �Mozӛ�?d!Y�B�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���~hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM9hjh))��}�(h,h/h0M9��h2h3h4hph<�h=Kub������       �                    �?� ��4d�?�           8�@              9                    �?��G�Vv�?.           �}@               8                    @.�ȓ�<�?U            �_@              +                    �?؇���X�?S            �]@                                   @xP�Fֺ�?>            @V@                                 �H@@4և���?'             L@                                   �?@9G��?!            �H@        ������������������������       �                     7@        	       
                 `f�)@$�q-�?             :@        ������������������������       �                     $@                                   �?      �?
             0@        ������������������������       �                     @                                   :@8�Z$���?	             *@        ������������������������       �                     �?                                  �*@�8��8��?             (@                                  B@      �?              @       ������������������������       �                     @                                   D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                    �?����X�?             @                                   K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �J@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?�'�`d�?            �@@       ������������������������       �                     4@               *                    ;@��
ц��?
             *@               )                   �8@      �?              @       !       "                 ���@���Q��?             @        ������������������������       �                     �?        #       (                   �6@      �?             @       $       '                 ��!@�q�q�?             @       %       &                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ,       7                    @z�G�z�?             >@       -       2                   �/@V�a�� �?             =@        .       /                     @      �?              @        ������������������������       �                      @        0       1                 ��'@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        3       6                 039@���N8�?             5@        4       5                 03�7@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     �?        ������������������������       �                      @        :       _                     �?1�}i��?�            �u@        ;       \                    �?؇>���?%            @P@       <       W                    �?��mo*�?"            �M@       =       D                    �?d,���O�?            �I@        >       ?                  Y>@r�q��?             (@        ������������������������       �                     �?        @       C                   �A@�C��2(�?             &@        A       B                 X�,@@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        E       R                   �J@�(�Tw��?            �C@       F       Q                   `@@���Q��?             9@       G       H                 �̌*@����X�?	             ,@        ������������������������       �                     �?        I       P                 �|�?@�θ�?             *@       J       K                    <@      �?             @        ������������������������       �                     �?        L       M                 �|Y=@���Q��?             @        ������������������������       �                     �?        N       O                 `fF<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        S       T                 `fF<@@4և���?             ,@        ������������������������       �                      @        U       V                   �Q@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        X       [                   �B@      �?              @        Y       Z                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ]       ^                  DdX@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        `       a                    $@��C���?�            �q@        ������������������������       �                      @        b       �                 �?�@h>#j�x�?�            �q@        c       �                   �@p��%���?S            @a@       d       e                     @���l��?>            �[@        ������������������������       �                     �?        f                        ��]@,�+�C�?=            �[@       g       ~                 �|�=@88��M�?:            �Z@       h       i                   �5@�m(�X�?-            @U@        ������������������������       �                     ,@        j       y                    �?h��@D��?%            �Q@       k       p                    �?�r����?            �F@        l       o                 ���@�t����?	             1@       m       n                   �7@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        q       t                 �|Y=@؇���X�?             <@        r       s                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        u       v                 ���@HP�s��?             9@        ������������������������       �                     @        w       x                 ��(@�����H�?
             2@       ������������������������       �      �?	             0@        ������������������������       �                      @        z       {                 �|�<@ ��WV�?             :@       ������������������������       �                     3@        |       }                 ��,@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     6@        �       �                   �:@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        �       �                   �C@^	����?_            @b@       �       �                     @@�0�!��?N            �]@        �       �                   �3@      �?             @@       �       �                   �)@؇���X�?             <@        �       �                    &@$�q-�?             *@       �       �                    5@ףp=
�?             $@        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|�<@z�G�z�?             .@        ������������������������       �                     @        �       �                 �|�=@�z�G��?             $@        ������������������������       �                      @        �       �                    @@      �?              @       ������������������������       �                     @        �       �                   �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|�=@�����?5            �U@       �       �                   �;@�LQ�1	�?*            @Q@       �       �                   �8@�<ݚ�?             B@       �       �                    �?��� ��?             ?@        ������������������������       �                     �?        �       �                 ��Y @�r����?             >@        �       �                 @3�@�q�q�?             (@        ������������������������       �                     @        �       �                    4@      �?              @       �       �                    1@�q�q�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             2@        �       �                 pf� @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 pf� @Pa�	�?            �@@        �       �                 �|Y=@$�q-�?	             *@        ������������������������       �                     �?        �       �                 ��) @�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     4@        �       �                   �@@X�<ݚ�?             2@       �       �                   �?@�q�q�?             "@        �       �                 �̌!@      �?             @       �       �                   �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��I @���Q��?             @        ������������������������       �                      @        �       �                 d�6@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 @3�@�<ݚ�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     ;@        �       �                     @`��
-��?�             m@        �       �                     �?d}h��?E             \@       �       �                    �?     ��?&             P@       �       �                    �?r�q��?             H@        �       �                    �?���N8�?             5@        ������������������������       �                     &@        �       �                    �?      �?             $@       �       �                 p"�X@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�����H�?             ;@       ������������������������       �        	             2@        �       �                 ��9L@�q�q�?             "@       �       �                 `�iJ@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?     ��?
             0@       �       �                    )@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                ����8@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             H@       �       �                    �?�C��2(�?             6@        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                   @B@�q�q�?             @       �       �                   �9@z�G�z�?             @        ������������������������       �                      @        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             .@        �       �                   �3@�θ�?             :@        �       �                 �z�'@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�KM�]�?             3@        ������������������������       �                     @        �       �                   �@@؇���X�?             ,@       �       �                    �?�8��8��?             (@        ������������������������       �                     @        �       �                    �?r�q��?             @       �       �                    1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    &@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       &                 ��8@dՔ���?J            @^@       �       �                 P�@b1<+�C�?-            @R@        ������������������������       �                     &@        �                          �?`՟�G��?'             O@        �                          �?�d�����?             3@       �       �                    �?�t����?	             1@       �       �                    �?�	j*D�?             *@       ������������������������       �                      @        �       �                 �|Y3@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?                                  �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                              03�1@��V#�?            �E@                               �/@�q�����?             9@                                �?     ��?             0@              
                P��%@և���X�?             @             	                  �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                              ��=)@�<ݚ�?             "@                                 �?�q�q�?             @                                7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �?�<ݚ�?             "@                               �0@���Q��?             @                             �|�:@      �?             @        ������������������������       �                     �?                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @              !                   �?�����H�?             2@                                 �?r�q��?             @        ������������������������       �                     �?                                 �3@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        "      #                ��i4@�8��8��?             (@        ������������������������       �                     @        $      %                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        '      8                   @�8��8��?             H@       (      /                   �?<���D�?            �@@        )      *                   �?���!pc�?	             &@        ������������������������       �                      @        +      ,                ��T?@�q�q�?             "@        ������������������������       �                     @        -      .                  @D@      �?             @        ������������������������       �                     @        ������������������������       �                     @        0      1                   @���7�?             6@        ������������������������       �                      @        2      7                ���A@P���Q�?             4@       3      4                   �?ףp=
�?             $@       ������������������������       �                      @        5      6                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     .@        �*       h�h))��}�(h,h/h0M9KK��h2h3h4hVh<�h=Kub��������������`uv��?,J>��?��VAm�?zR}%��?M&��d2�?m6��f��?�$I�$I�?۶m۶m�?�я~���?�.p��?�$I�$I�?n۶m۶�?9/���?������?              �?;�;��?�؉�؉�?              �?      �?      �?              �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?      �?                      �?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?        '�l��&�?6�d�M6�?              �?�;�;�?�؉�؉�?      �?      �?�������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?                      �?      �?        �������?�������?a���{�?��{a�?      �?      �?              �?�������?UUUUUU�?              �?      �?        �a�a�?��y��y�?      �?      �?              �?      �?                      �?              �?      �?        q�a���?<y�#�?�����? �����?�<�"h�?W'u_�?�������?PPPPPP�?�������?UUUUUU�?              �?]t�E�?F]t�E�?�������?�������?      �?                      �?      �?        �o��o��?� � �?333333�?�������?�$I�$I�?�m۶m��?      �?        �؉�؉�?ى�؉��?      �?      �?              �?333333�?�������?      �?              �?      �?      �?                      �?              �?      �?        n۶m۶�?�$I�$I�?      �?        �������?UUUUUU�?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��YR��?��3m���?              �?p�z2~��?�D+l$�?�g��%�?ہ�v`��?��蕱�?5'��Ps�?      �?        �}��7��?��)A��?+J�#��?����f��?]]]]]]�?�?      �?        ��V��?�'�K=�?�������?�?<<<<<<�?�?      �?      �?              �?      �?              �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?q=
ףp�?{�G�z�?      �?        �q�q�?�q�q�?      �?      �?      �?        O��N���?;�;��?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        [�lٲe�?�&M�4i�?ZZZZZZ�?�������?      �?      �?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?�������?�������?      �?      �?      �?              �?        �������?�������?      �?        ffffff�?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ;���C��?/�I��?��Moz��?Y�B��?9��8���?�q�q�?�{����?�B!��?      �?        �������?�?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?      �?                      �?|���?|���?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        r�q��?�q�q�?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?                      �?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?              �?        ����S��?Ⱥ��X��?�$I�$I�?�m۶m��?      �?     ��?UUUUUU�?�������?��y��y�?�a�a�?              �?      �?      �?      �?      �?              �?      �?              �?        �q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?F]t�E�?]t�E�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?ى�؉��?�؉�؉�?۶m۶m�?�$I�$I�?              �?      �?        �k(���?(�����?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?              �?      �?        ��J���?���k���?�;w�ܹ�?Ĉ#F��?      �?        �1�c��?�s�9��?y�5���?Cy�5��?�������?�������?;�;��?vb'vb'�?              �?�������?�������?      �?                      �?      �?      �?              �?      �?                      �?eMYS֔�?6eMYS��?�p=
ף�?���Q��?      �?      �?�$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        �q�q�?9��8���?�������?333333�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�q�q�?�q�q�?�������?UUUUUU�?      �?        �������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?|���?|���?F]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �.�袋�?F]t�E�?      �?        ffffff�?�������?�������?�������?      �?              �?      �?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJCLUhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                     @�t����?�           8�@               7                   �<@�h��?�             t@                                   :@Dc}h���?<             \@                                   �?�5��?             K@                                 �;@X�<ݚ�?             B@                                  �?     ��?             @@                                 �2@R�}e�.�?             :@        ������������������������       �                     @        	                           �?��Q��?             4@        
                        pf�,@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @                                  �'@���!pc�?	             &@                                   �?���Q��?             @        ������������������������       �                      @                                  �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?�����H�?             2@        ������������������������       �                     &@                                   ,@����X�?             @       ������������������������       �                     @        ������������������������       �                      @               ,                    �?�y��*�?!             M@              )                 ��X@��(\���?             D@              (                    �?XB���?             =@               !                    �?���N8�?             5@       ������������������������       �                     (@        "       #                    �?�����H�?             "@        ������������������������       �                      @        $       %                   �;@؇���X�?             @        ������������������������       �                      @        &       '                 `f�D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        *       +                    �?"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        -       0                    �?�<ݚ�?             2@       .       /                  "&d@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        1       6                    �?      �?              @       2       5                     �?r�q��?             @       3       4                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        8       �                    �?\qr��?�            @j@       9       j                     �?V{q֛w�?s            @g@       :       [                    �?���0��?C             [@       ;       @                    �?l�;�	�?-            �R@        <       ?                 �iE@��S�ۿ?
             .@        =       >                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        A       L                    �?��0u���?#             N@        B       C                   @@@���y4F�?
             3@        ������������������������       �                     "@        D       K                 @�Cq@���Q��?             $@       E       F                 `v�<@      �?              @        ������������������������       �                     �?        G       J                 p�i@@؇���X�?             @        H       I                    H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        M       Z                   �Q@�4F����?            �D@       N       Y                  )?@�(�Tw��?            �C@       O       P                 �|Y=@��>4և�?             <@        ������������������������       �                     @        Q       R                 03:@r�q��?             8@        ������������������������       �                     @        S       X                   @=@ҳ�wY;�?
             1@       T       W                 `f�;@��
ц��?	             *@       U       V                   �J@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             &@        ������������������������       �                      @        \       ]                    �?���!pc�?            �@@       ������������������������       �                     2@        ^       a                    �?���Q��?	             .@        _       `                   �H@      �?             @        ������������������������       �                      @        ������������������������       �                      @        b       c                  x#J@���|���?             &@        ������������������������       �                     @        d       e                    A@      �?              @        ������������������������       �                      @        f       g                   �B@�q�q�?             @        ������������������������       �                      @        h       i                   �E@      �?             @        ������������������������       �                      @        ������������������������       �                      @        k       �                   �E@�q�q�?0            �S@       l       {                    �?�f7�z�?$             M@       m       p                 �|�=@�>$�*��?            �D@        n       o                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        q       x                   �A@�'�=z��?            �@@       r       s                    �?�q�q�?             2@        ������������������������       �                      @        t       w                    @@      �?
             0@       u       v                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        y       z                    �?�q�q�?             .@        ������������������������       �                     @        ������������������������       �                     $@        |       }                    �?ҳ�wY;�?             1@        ������������������������       �                     @        ~                          �7@      �?             (@        ������������������������       �                     �?        �       �                   �?@�eP*L��?             &@        ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?ףp=
�?             4@        �       �                    5@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             0@        �       �                    �?�q�q�?             8@       ������������������������       �                     0@        ������������������������       �                      @        �       �                    /@��VI��?�            Px@        �       �                    @*O���?             B@       �       �                    @8�Z$���?             :@       ������������������������       �        	             ,@        �       �                 �&�)@�q�q�?             (@        ������������������������       �                     @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?ףp=
�?	             $@        ������������������������       �                     @        �       �                    @z�G�z�?             @        ������������������������       �                      @        �       �                 ��T?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�]�5�?�            v@        �       �                    �?�eP*L��?;            �X@        �       �                    �?z�G�z�?            �F@       �       �                    �?���"͏�?            �B@        �       �                 �|Y=@�q�q�?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�חF�P�?             ?@       �       �                 �|�9@@4և���?             <@        ������������������������       �                     $@        �       �                  ��@�����H�?             2@        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?r�q��?%             K@       �       �                 �|Y=@      �?              H@        �       �                    5@      �?              @        �       �                 �{@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @       �       �                   �6@      �?             @        ������������������������       �                      @        �       �                 xF*@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�=@�(\����?             D@       �       �                 ���@XB���?             =@        �       �                    �?$�q-�?	             *@       �       �                 ���@�����H�?             "@       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     0@        ������������������������       �                     &@        �       �                 �|Y7@      �?             @        ������������������������       �                     �?        �       �                    �?���Q��?             @        �       �                 ��.@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                  �v6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @Q!@J�:�Ȣ�?�            �o@       �       �                    �?�K�	H�?\             c@       �       �                    �?�T�2�?[            �b@        �       �                    ;@��.k���?             1@       �       �                   �6@z�G�z�?             $@        ������������������������       �                     @        �       �                   �9@�q�q�?             @       �       �                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?����e��?P            �`@       �       �                 ��) @�-.�1a�?J            �^@       �       �                   �0@@m���?E             ]@        �       �                 pf�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        C            @\@        �       �                 �|Y8@؇���X�?             @        ������������������������       �                     @        �       �                 ��y @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        �                         @B@N��>��?C            @Y@       �                       �|�=@̠�4��?6            �T@       �                       ��Y1@�'�`d�?+            �P@       �                          �?��i#[�?             E@       �       �                    �?��Q���?             D@       �       �                 @3�!@������?             A@        �       �                    �?և���X�?             @       �       �                    6@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 @33/@PN��T'�?             ;@       �       �                   �2@�}�+r��?             3@        �       �                 �yW#@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        �       �                 �|�;@      �?              @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �#@      �?             @        ������������������������       �                     �?        �                           �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                 �? �q�q�?             8@        ������������������������       �                     $@              
                   ;@@4և���?	             ,@             	                   �?؇���X�?             @                                 9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                              �T)D@ҳ�wY;�?             1@                               �*@և���X�?
             ,@                                 @@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                �A@X�<ݚ�?             "@                               @.@      �?              @        ������������������������       �                      @                                �>@      �?             @        ������������������������       �                     �?                                  @���Q��?             @                                �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������G�+J>�?r%�k���?�.>9�?��h�`��?%I�$I��?n۶m۶�?/�����?h/�����?r�q��?�q�q�?      �?      �?'vb'vb�?�;�;�?      �?        �������?ffffff�?r�q��?�q�q�?              �?      �?        F]t�E�?t�E]t�?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?              �?      �?        �q�q�?�q�q�?              �?�$I�$I�?�m۶m��?              �?      �?        GX�i��?�4�rO#�?333333�?�������?�{a���?GX�i���?�a�a�?��y��y�?              �?�q�q�?�q�q�?              �?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?                      �?F]t�E�?/�袋.�?              �?      �?        �q�q�?9��8���?333333�?ffffff�?              �?      �?              �?      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�8�8�?�؏�؏�?B!��?�{����?���Kh�?����K�?ƒ_,���?t�@�t�?�?�������?      �?      �?      �?                      �?              �?�������?""""""�?6��P^C�?(������?      �?        333333�?�������?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?ە�]���?KԮD�J�?�o��o��?� � �?۶m۶m�?I�$I�$�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?�؉�؉�?�;�;�?F]t�E�?]t�E]�?              �?      �?              �?                      �?      �?                      �?t�E]t�?F]t�E�?              �?333333�?�������?      �?      �?              �?      �?        ]t�E]�?F]t�E�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?O#,�4��?a���{�?�18���?�����?      �?      �?              �?      �?        |���?|��|�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?              �?      �?      �?        ]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?              �?      �?        �������?�������?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        ���k�2�?}�$(���?�q�q�?�q�q�?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?�������?�������?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?zXF��b�?��|u�?t�E]t�?]t�E�?�������?�������?*�Y7�"�?v�)�Y7�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��RJ)��?�Zk����?�$I�$I�?n۶m۶�?              �?�q�q�?�q�q�?      �?                      �?      �?                      �?�������?UUUUUU�?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?      �?              �?      �?      �?      �?                      �?              �?333333�?�������?GX�i���?�{a���?�؉�؉�?;�;��?�q�q�?�q�q�?      �?              �?      �?      �?              �?              �?              �?      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?�b�X,�?�t:�N��?�g�g�?�l�l�?��*�3��?7`��c.�?�������?�?�������?�������?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �>����?|���?{����z�?�h
���?�{a��?�{a���?UUUUUU�?UUUUUU�?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�be�F�?�tj��?�����\�?]V��F�?6�d�M6�?'�l��&�?�a�a�?�<��<��?333333�?�������?xxxxxx�?�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        &���^B�?h/�����?�5��P�?(�����?      �?      �?      �?                      �?      �?              �?      �?      �?              �?      �?              �?      �?              �?      �?              �?333333�?�������?              �?      �?                      �?�������?UUUUUU�?      �?        n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?۶m۶m�?�$I�$I�?�������?�������?              �?      �?        r�q��?�q�q�?      �?      �?      �?              �?      �?      �?        �������?333333�?      �?      �?              �?      �?                      �?              �?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������                           @S*f���?�           8�@                                @3�4@�<ݚ�?            �F@        ������������������������       �        
             0@                                   �?J�8���?             =@                                   �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   @      �?             8@       	                            @�����?             3@       
                           �?�8��8��?             (@       ������������������������       �                     "@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                ��T?@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                  @�bI����?�           Є@                                @L@ k��p2�?�           h�@              r                    �?����?�           Ѓ@               W                 �DhF@"��z��?w            �g@              &                 ���@O����?U             b@               %                    �?�?�'�@�?             C@              $                    �?r�q��?             >@                                  �?�+$�jP�?             ;@        ������������������������       �                     �?               !                 ���@8�Z$���?             :@                                  �7@�C��2(�?             &@                                   5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        "       #                 �|=@z�G�z�?             .@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        '       P                    �?��k��?A            �Z@       (       E                    �?��
ц��?7            �V@       )       6                     @�^�����?'             O@        *       -                    �?�ՙ/�?             5@        +       ,                     �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        .       5                    C@      �?             ,@       /       2                 ���<@�z�G��?             $@       0       1                   @@@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        3       4                 ��tA@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        7       D                 �|Y?@�p ��?            �D@       8       9                    �?      �?             @@       ������������������������       �                     2@        :       ?                 �|�;@؇���X�?
             ,@        ;       <                 �y�*@�q�q�?             @        ������������������������       �                     �?        =       >                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        @       C                 ��(@�C��2(�?             &@       A       B                 ���@      �?              @        ������������������������       �                      @        ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �                     "@        F       K                    �?8^s]e�?             =@        G       J                   �-@�����H�?             "@        H       I                   �,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        L       M                  �v6@P���Q�?	             4@       ������������������������       �                     *@        N       O                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        Q       R                     @���Q��?
             .@        ������������������������       �                     @        S       V                    �?���Q��?             $@       T       U                    3@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        X       c                 �UcV@�㙢�c�?"             G@        Y       Z                 p�1N@�8��8��?             8@        ������������������������       �                      @        [       `                    �?      �?             0@       \       _                   �9@$�q-�?
             *@        ]       ^                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        a       b                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        d       e                    �?���!pc�?             6@        ������������������������       �        	             (@        f       g                   �1@���Q��?	             $@        ������������������������       �                      @        h       q                    D@      �?              @       i       n                    �?���Q��?             @       j       m                    �?�q�q�?             @       k       l                 �̾w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        o       p                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        s       �                    �?<=�h)W�?           �{@        t       �                  �#@�Kǔ�{�?a            `d@        u       z                   �@      �?             @@        v       y                 ��@؇���X�?             ,@       w       x                 �|Y:@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        {       �                    �?�<ݚ�?             2@       |       �                  SE"@@�0�!��?
             1@       }       �                 ��� @      �?              @       ~       �                    �?����X�?             @              �                 �?�@���Q��?             @        ������������������������       �                     �?        �       �                   �8@      �?             @        ������������������������       �                     �?        �       �                 �|�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?D����\�?O            ``@       �       �                     @�~i��?@            @[@       �       �                     �?x��B�R�?2            �V@        ������������������������       �                     :@        �       �                    �?P�2E��?$            @P@       �       �                   �;@��<D�m�?            �H@        �       �                   �5@z�G�z�?             $@        ������������������������       �                     @        �       �                    �?����X�?             @        �       �                   �'@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �E@ ���J��?            �C@       ������������������������       �                     ?@        �       �                   @F@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             0@        �       �                   �D@      �?             2@       �       �                    �?     ��?             0@       �       �                 03�1@�z�G��?             $@       �       �                 �|�;@�<ݚ�?             "@        �       �                    4@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        �       �                    1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `fv1@      �?             @        ������������������������       �                      @        �       �                 `fV6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���|���?             6@        �       �                 ���0@      �?             @        ������������������������       �                      @        �       �                      @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @�E��ӭ�?             2@        ������������������������       �                     @        ������������������������       �        	             *@        �       �                 ��$:@hk��E�?�            �q@       �       �                 ��@0�%�J�?�            �k@        ������������������������       �                     D@        �       �                   �<@�D����?s            �f@        �       �                    �?�k~X��?0             R@       �       �                     @ _�@�Y�?'             M@        ������������������������       �                      @        �       �                   �2@p���?!             I@        �       �                   �1@      �?              @        ������������������������       �                     @        �       �                 ��@z�G�z�?             @        ������������������������       �                     @        �       �                 ��Y @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     E@        ������������������������       �        	             ,@        �       �                   �?@�:�H:�?C            @[@        �       �                    �?�>4և��?              L@       �       �                     @r�����?            �J@        �       �                   �'@�����H�?             "@        ������������������������       �                     @        �       �                     �?z�G�z�?             @        ������������������������       �                     �?        �       �                 �|�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �>@�������?             F@       �       �                 ��L@�S����?             C@        ������������������������       �      �?             @        �       �                 �|Y=@     ��?             @@        �       �                 ���"@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�=@@4և���?             <@       �       �                 ��) @���7�?             6@       ������������������������       �                     ,@        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �̌!@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 pff@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �D@�O4R���?#            �J@       ������������������������       �                    �A@        �       �                   @E@�X�<ݺ?             2@        �       �                     @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             .@        �                           �?�q�q�?&             N@       �                         �J@      �?             G@       �       
                  �G@�>$�*��?            �D@       �       �                 �T!@@��.k���?             A@        �       �                 �|�<@z�G�z�?             $@        ������������������������       �                     @        �       �                 X�,@@����X�?             @        �       �                 `fF<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 03k:@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        �       	                03�U@�q�q�?             8@       �                       ��yC@���N8�?             5@                                 �A@      �?             @       ������������������������       �                     @        ������������������������       �                     @                              �|Y>@�r����?
             .@        ������������������������       �                     @                                 A@�<ݚ�?             "@                                @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                �7@؇���X�?
             ,@        ������������������������       �                     @                              0�E@      �?              @        ������������������������       �                      @                                 ;@�q�q�?             @        ������������������������       �                     �?                              �|�>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     *@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������H�7�?=�o�a��?�q�q�?9��8���?              �?|a���?�rO#,��?�������?�������?      �?                      �?      �?      �?^Cy�5�?Q^Cy��?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�m۶m��?�$I�$I�?      �?                      �?              �?�@\�9	�?�~G����?�cEK@��?8uig�?�C!�n�?Txǽ�"�?�
��v��?q�����?��8��8�?�8��8��?������?y�5���?�������?UUUUUU�?/�����?B{	�%��?              �?;�;��?;�;��?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?        �������?�������?      �?              �?      �?      �?              �?        oe�Cj��?"5�x+��?�;�;�?�؉�؉�?���{��?!�B�?�a�a�?�<��<��?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?ffffff�?333333�?۶m۶m�?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?dp>�c�?8��18�?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?]t�E�?F]t�E�?      �?      �?      �?        �������?UUUUUU�?      �?              �?        |a���?	�=����?�q�q�?�q�q�?      �?      �?              �?      �?                      �?ffffff�?�������?      �?        ۶m۶m�?�$I�$I�?      �?                      �?333333�?�������?      �?        �������?333333�?      �?      �?      �?                      �?      �?        d!Y�B�?�7��Mo�?UUUUUU�?UUUUUU�?              �?      �?      �?;�;��?�؉�؉�?UUUUUU�?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        t�E]t�?F]t�E�?              �?333333�?�������?              �?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?      �?        �I .Ԝ�?el��W��?kq�}�?�uǋ-��?      �?      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?9��8���?�q�q�?ZZZZZZ�?�������?      �?      �?�m۶m��?�$I�$I�?333333�?�������?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?                      �?�U���g�?���[��?��A��.�?��w� z�?��?�����?              �?z�z��?_�^��?և���X�?��S�r
�?�������?�������?              �?�$I�$I�?�m۶m��?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �A�A�?��-��-�?              �?      �?      �?      �?                      �?              �?      �?      �?      �?      �?333333�?ffffff�?�q�q�?9��8���?      �?      �?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?              �?        ]t�E]�?F]t�E�?      �?      �?              �?      �?      �?              �?      �?        �q�q�?r�q��?              �?      �?        ՆL�V��?���Υ��?~/C~/C�?�ͫ?      �?        B-`L���?������?�8��8��?�q�q�?#,�4�r�?�{a���?      �?        \���(\�?{�G�z�?      �?      �?      �?        �������?�������?      �?              �?      �?              �?      �?              �?              �?        Ṷ�H��?\����չ?�$I�$I�?�m۶m��?Dj��V��?�V�9�&�?�q�q�?�q�q�?      �?        �������?�������?      �?              �?      �?              �?      �?        t�E]t�?/�袋.�?(������?^Cy�5�?      �?      �?      �?      �?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?�.�袋�?F]t�E�?      �?              �?      �?              �?      �?        �������?UUUUUU�?      �?                      �?      �?      �?      �?                      �?      �?        :�&oe�?�x+�R�?      �?        ��8��8�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?      �?      �?�����?�18���?�������?�?�������?�������?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?�a�a�?��y��y�?      �?      �?      �?                      �?�������?�?      �?        9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ"�a,hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������       
                    @�����?�           8�@                                    @���B���?"             J@        ������������������������       �                     9@                                   @��}*_��?             ;@        ������������������������       �        
             *@                                ��T?@����X�?
             ,@       ������������������������       �                      @               	                 ���A@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @               `                    �?�oH'0��?�           ��@               )                     @ �o_��?�             l@              (                    �? d�=��?O            @\@              '                 0Cd=@�Zl�i��?7            @T@                                  �B@z�G�z�?             D@                                 �;@�>����?             ;@                                   �?"pc�
�?             &@        ������������������������       �                     @                                  �'@�q�q�?             @        ������������������������       �                     @                                  �9@�q�q�?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@               "                  ��9@��
ц��?             *@              !                   �,@�q�q�?             "@                                  �'@      �?             @                                 �J@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        #       &                    �?      �?             @       $       %                    K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �D@        ������������������������       �                     @@        *       +                    )@ �Cc��?F             \@        ������������������������       �                     @        ,       S                    �?�xGZ���?B            @Z@       -       8                  ��@L�qA��?/            �R@        .       /                    8@\-��p�?             =@        ������������������������       �                     "@        0       5                    �?z�G�z�?             4@       1       4                  ��@�t����?	             1@        2       3                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        6       7                 �&B@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        9       F                 �|�;@
;&����?             G@        :       ?                    �?      �?             8@        ;       <                 �&�)@����X�?             @        ������������������������       �                     @        =       >                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        @       A                  �#@�IєX�?
             1@       ������������������������       �                     &@        B       E                    �?r�q��?             @        C       D                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        G       N                    �?���!pc�?             6@        H       M                   &@և���X�?             @       I       J                 ��� @z�G�z�?             @        ������������������������       �                      @        K       L                    A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        O       P                 �|Y>@�r����?
             .@       ������������������������       �                     &@        Q       R                    @@      �?             @        ������������������������       �                      @        ������������������������       �                      @        T       _                 ���7@�q�q�?             >@       U       Z                    �?j���� �?             1@        V       Y                    �?      �?              @       W       X                 `�@1@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        [       \                   �;@�����H�?             "@       ������������������������       �                     @        ]       ^                   �=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        a       �                     �?\����?            {@        b       g                   �<@P��MO�?5            �T@        c       d                   �8@���!pc�?             &@        ������������������������       �                      @        e       f                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        h       �                 p�w@�<ݚ�?-             R@       i       v                    �?z�G�z�?,            �Q@        j       s                    �?"pc�
�?             6@       k       r                 ��2>@      �?
             0@        l       m                 ���<@�����H�?             "@        ������������������������       �                     @        n       q                    �?      �?             @       o       p                 X��E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        t       u                 @�pX@      �?             @       ������������������������       �                     @        ������������������������       �                     @        w       �                    �?�q�q�?             H@       x       �                   �>@��k=.��?            �G@       y       �                   @>@�q�q�?             ;@       z       {                 03:@      �?             8@        ������������������������       �                     @        |       �                    R@�z�G��?             4@       }       ~                 03k:@�d�����?             3@        ������������������������       �                     �?               �                    J@�<ݚ�?
             2@       �       �                 `f�;@�q�q�?             (@       �       �                   @G@      �?              @       �       �                   �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �z�G�z�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?TO$�?�            �u@       �       �                     @�luL3�?�            Ps@        �       �                    4@Pa�	�?)            �P@        �       �                   �2@؇���X�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                   �@@P����?%            �M@       ������������������������       �                     A@        �       �                   �*@`2U0*��?             9@       �       �                   �)@��S�ۿ?	             .@        ������������������������       �                     "@        �       �                   �A@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     $@        �       �                 �T)D@��L9���?�            `n@       �       �                    �?�*/�8V�?�            `m@        �       �                 �|Y=@����X�?             5@        �       �                    �?�q�q�?             "@       �       �                    ;@      �?              @       �       �                   �7@���Q��?             @       �       �                    5@      �?             @       �       �                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             (@        �       �                 0SE @p7Y���?�            �j@       �       �                    �?���C��?g            �c@        �       �                 �|Y=@r�q��?             8@        ������������������������       �                      @        �       �                 �Y�@�C��2(�?             6@        ������������������������       �                     @        �       �                 ��(@�t����?             1@       �       �                 X��A@      �?
             0@       ������������������������       �8�Z$���?             *@        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��) @�Aʑ���?X            �`@       �       �                   @4@ՀJ��?W            �`@        �       �                   �2@����X�?             5@        �       �                 pf�@      �?              @        ������������������������       �                     @        �       �                    1@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        �       �                    �?�θ�?	             *@       �       �                 @3�@r�q��?             (@       ������������������������       �                      @        �       �                   �3@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �8@�h����?H             \@        �       �                    �?ȵHPS!�?             :@       �       �                    7@�LQ�1	�?             7@       ������������������������       �        
             .@        �       �                 `fF@      �?              @        �       �                 �&b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �>@��+��<�?9            �U@       ������������������������       �        !            �I@        �       �                   �?@�#-���?            �A@        ������������������������       �                      @        �       �                 �?�@Pa�	�?            �@@       ������������������������       �                     7@        �       �                   �@@ףp=
�?             $@        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���!@ �Jj�G�?%            �K@        �       �                 @Q!@�IєX�?             1@        ������������������������       �                      @        �       �                    8@��S�ۿ?	             .@       ������������������������       �                     $@        �       �                 �|Y<@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     C@        �       �                    ;@      �?              @        ������������������������       �                     @        �       �                 �|�>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|Y>@؇���X�?             E@       �       �                 �̌4@�<ݚ�?             ;@        �       �                 ��*@և���X�?             ,@        ������������������������       �                     @        �       �                    �?�q�q�?             "@        ������������������������       �                      @        �       �                 8#�1@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �        
             .@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub������������������?��܍��?ى�؉��?��؉���?              �?B{	�%��?_B{	�%�?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        /X���+�?�O��4��?�Q����?
ףp=
�?x�!���?���	��?�����H�?�"e����?�������?�������?h/�����?�Kh/��?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?�؉�؉�?�;�;�?UUUUUU�?UUUUUU�?      �?      �?�������?333333�?              �?      �?              �?                      �?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?        �A�A�?�_�_�?�K~���?t�@��?�{a���?a����?              �?�������?�������?�?<<<<<<�?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?Y�B��?�Mozӛ�?      �?      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?�?�?      �?        �������?UUUUUU�?      �?      �?              �?      �?              �?        t�E]t�?F]t�E�?�$I�$I�?۶m۶m�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�?�������?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?ZZZZZZ�?�������?      �?      �?۶m۶m�?�$I�$I�?      �?                      �?              �?�q�q�?�q�q�?              �?      �?      �?      �?                      �?      �?        \.���?��G����?��7�:��?���ˊ��?t�E]t�?F]t�E�?      �?        �q�q�?�q�q�?              �?      �?        9��8���?�q�q�?�������?�������?/�袋.�?F]t�E�?      �?      �?�q�q�?�q�q�?      �?              �?      �?      �?      �?              �?      �?              �?              �?              �?      �?              �?      �?        UUUUUU�?�������?g���Q��?br1���?UUUUUU�?UUUUUU�?      �?      �?      �?        ffffff�?333333�?Cy�5��?y�5���?              �?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?              �?                      �?              �?      �?                      �?              �?���t��?ƯQpZ��?�+&��?NZ�Ϯ�?|���?|���?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?�V'u�?'u_[�?      �?        ���Q��?{�G�z�?�������?�?      �?        �������?UUUUUU�?      �?      �?      �?              �?        �ϙZ.�?﯃1+��?r1����?m�w6�;�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?�������?333333�?      �?      �?      �?      �?      �?                      �?              �?      �?                      �?      �?              �?        ���B�(�?�#蝺�?\�琚`�?"5�x+��?�������?UUUUUU�?              �?]t�E�?F]t�E�?      �?        <<<<<<�?�?      �?      �?;�;��?;�;��?      �?              �?        ���u��?Ũ�oS��?��7G��?�qA��?�m۶m��?�$I�$I�?      �?      �?      �?              �?      �?      �?      �?              �?ى�؉��?�؉�؉�?�������?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?��N��N�?�؉�؉�?��Moz��?Y�B��?      �?              �?      �?      �?      �?      �?                      �?      �?              �?        �#�;��?w�qGܡ?      �?        �A�A�?_�_�?              �?|���?|���?      �?        �������?�������?�������?�������?      �?                      �?k߰�k�?��)A��?�?�?      �?        �������?�?      �?        �������?�������?              �?      �?              �?              �?      �?              �?�������?�������?      �?                      �?۶m۶m�?�$I�$I�?9��8���?�q�q�?�$I�$I�?۶m۶m�?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�8�hhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM=hjh))��}�(h,h/h0M=��h2h3h4hph<�h=Kub������       �                     @��t���?�           8�@               y                  x#J@����>��?�            ps@              j                    �?T�$@��?�            �j@              /                   �2@�t���?l            �e@                                   @�f���?2            �T@        ������������������������       �                      @               .                    �?�EH,���?,            �R@              -                    L@��+��?+            �R@       	       &                   �C@��.k���?&             Q@       
                           &@�>���?             K@                                  �5@8�A�0��?	             6@                                   �?"pc�
�?             &@        ������������������������       �                     @        ������������������������       �����X�?             @                                   �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @                                  �;@      �?             @@        ������������������������       �                     (@                                   �?���Q��?             4@        ������������������������       �                     �?                                   �?p�ݯ��?             3@        ������������������������       �                     �?                                  @@@b�2�tk�?             2@                                   �?r�q��?             @       ������������������������       �                     @                                �|�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                `fF)@      �?             (@        ������������������������       �                      @                #                    �?���Q��?             $@        !       "                   �B@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        $       %                   �A@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        '       ,                   �*@d}h���?             ,@       (       )                    �?      �?              @        ������������������������       �                     @        *       +                   �F@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        0       5                   �9@�μ���?:            @V@        1       2                     �?z�G�z�?             @        ������������������������       �                      @        3       4                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        6       c                    H@d}h���?6             U@       7       F                 �|Y=@�㙢�c�?+            @Q@        8       ?                    �?X�Cc�?	             ,@        9       >                     �?����X�?             @       :       ;                   @>@      �?             @        ������������������������       �                     �?        <       =                 `ffC@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        @       A                    <@և���X�?             @        ������������������������       �                     �?        B       C                   �7@      �?             @        ������������������������       �                      @        D       E                 0C�:@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        G       b                   �F@X�;�^o�?"            �K@       H       S                    �?���V��?            �F@        I       J                 �|�=@�<ݚ�?             "@        ������������������������       �                     @        K       R                   �A@���Q��?             @       L       Q                    �?      �?             @       M       N                 `f&;@�q�q�?             @        ������������������������       �                     �?        O       P                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        T       a                   @F@4?,R��?             B@       U       Z                    �?�t����?             A@        V       Y                   �C@���Q��?             @       W       X                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        [       `                     �?XB���?             =@       \       _                 �̤<@�IєX�?             1@        ]       ^                 X�,@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     (@        ������������������������       �      �?              @        ������������������������       �                     $@        d       e                    �?���Q��?             .@        ������������������������       �                     @        f       g                   �J@"pc�
�?	             &@        ������������������������       �                     �?        h       i                   �R@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        k       l                    �?(L���?            �E@       ������������������������       �                     <@        m       n                     �?���Q��?             .@        ������������������������       �                     �?        o       p                   `6@X�Cc�?
             ,@        ������������������������       �                     @        q       t                 �D0@@�eP*L��?             &@       r       s                    1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        u       x                    �?z�G�z�?             @       v       w                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        z       �                    �?�q�Q�?=             X@        {       �                     �?�X����?             F@       |       �                    �?�^�����?            �E@       }       ~                    �?����"�?             =@       ������������������������       �        
             .@               �                 �\@d}h���?             ,@        �       �                 03/O@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �       �                 �|�9@؇���X�?
             ,@        ������������������������       �                     @        �       �                  �k@�<ݚ�?             "@       �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?4��?�?              J@       ������������������������       �                     ?@        �       �                   �H@���N8�?             5@       �       �                    A@      �?
             0@        ������������������������       �                      @        �       �                 `ށK@      �?              @        �       �                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `f^@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       <                   @�+e�X�?�             y@       �       �                    �?LZ���?�            px@        �       �                    �?N{�T6�?F            �[@        �       �                    �?���� �?            �D@        �       �                 P��+@և���X�?             5@        ������������������������       �                     @        �       �                    �?     ��?             0@        �       �                 ���,@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Q��?             $@       �       �                 83�0@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y=@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 X�,A@ףp=
�?             4@       �       �                    �?�}�+r��?             3@       �       �                 �|Y8@@4և���?	             ,@        ������������������������       �                     @        �       �                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 P�J@�㙢�c�?.            @Q@       �       �                    �?ףp=
�?             D@        �       �                   �6@؇���X�?
             ,@        �       �                 �{@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        �       �                  ��@$�q-�?             :@        ������������������������       �                     "@        �       �                 �|Y=@�t����?             1@        ������������������������       �                     �?        �       �                 X��A@      �?             0@       ������������������������       ���S�ۿ?
             .@        ������������������������       �                     �?        �       �                 03�7@�c�Α�?             =@       �       �                 =
�@���|���?             6@        ������������������������       �                      @        �       �                    �?�z�G��?             4@       �       �                   �;@@�0�!��?             1@        ������������������������       �                     @        �       �                  �v6@�θ�?
             *@       �       �                 �|Y=@�C��2(�?	             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��}@hX͇���?�            �q@        ������������������������       �                     A@        �                       ���"@�����?�            �n@       �       �                    �?     ��?Z             b@        �       �                    �?�G�z��?             4@       �       �                 @3�@D�n�3�?             3@       �       �                    ;@և���X�?
             ,@       �       �                    �?z�G�z�?             $@       �       �                   �9@�<ݚ�?             "@       �       �                   �7@      �?             @       �       �                 P��@�q�q�?             @        ������������������������       �                     �?        �       �                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �                          �?���-T��?M             _@       �       �                 �?�@����n�?I            �]@        �       �                   �@dP-���?            �G@       �       �                 �|�<@�r����?             >@       ������������������������       �                     3@        �       �                   @@@���|���?             &@       �       �                 �&B@      �?              @       �       �                 �|Y>@�q�q�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     1@        �                       ���!@tk~X��?*             R@       �       �                 �|Y<@��a�n`�?%             O@        �       �                   �9@
j*D>�?             :@       �       �                 0S5 @�X����?             6@       �       �                   �3@     ��?
             0@        �       �                    1@�z�G��?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �                        @3�@�8��8��?             B@        �       �                   �?@�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �A@      �?              @        ������������������������       �                     @        ������������������������       ��q�q�?             @                              ��) @ 7���B�?             ;@       ������������������������       �                     7@                              ��y @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @              3                �|�=@�ެD��?D            �Y@       	                         @�Y�����?7            �T@        
                      ���A@�q�q�?
             (@                             ��T?@�z�G��?             $@                                 @      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @              &                   �?D��\��?-            �Q@                                 #@r٣����?            �@@        ������������������������       �                     �?                                �#@     ��?             @@                                �<@�q�q�?             (@                                �?      �?              @                                 4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                              �|Y=@      �?             @        ������������������������       �                     @        ������������������������       �                     �?              #                   �?R���Q�?             4@             "                   ;@      �?
             0@               !                �!&B@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        $      %                ��l4@      �?             @        ������������������������       �                      @        ������������������������       �                      @        '      2                   �?�}�+r��?             C@        (      -                   �?�KM�]�?             3@       )      ,                   �?@4և���?             ,@        *      +                �|�;@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        .      1                   �?z�G�z�?             @        /      0                   +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        4      5                0S�*@      �?             4@        ������������������������       �                     @        6      ;                   @����X�?             ,@       7      :                   �?r�q��?
             (@        8      9                  �B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        �*       h�h))��}�(h,h/h0M=KK��h2h3h4hVh<�h=Kub�������������nԾ���?5"W��6�?��f�?t�����?�b?-��?X:Ɂ���?A_���?}A_���?"�%��?�������?      �?        7�i�6�?�_,�Œ�?�S�n�?*�Y7�"�?�?�������?��Kh/�?�Kh/��?/�袋.�?颋.���?F]t�E�?/�袋.�?              �?�$I�$I�?�m۶m��?]t�E]�?F]t�E�?              �?      �?              �?      �?      �?        �������?333333�?      �?        Cy�5��?^Cy�5�?              �?9��8���?�8��8��?UUUUUU�?�������?              �?      �?      �?              �?      �?              �?      �?      �?        �������?333333�?UUUUUU�?�������?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?I�$I�$�?      �?      �?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�\��?�я~���?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        I�$I�$�?۶m۶m�?�7��Mo�?d!Y�B�?%I�$I��?�m۶m��?�m۶m��?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �$I�$I�?۶m۶m�?      �?              �?      �?      �?              �?      �?              �?      �?        �־a��?J��yJ�?[�[��?�>�>��?9��8���?�q�q�?      �?        333333�?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?              �?        �8��8��?r�q��?<<<<<<�?�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?GX�i���?�{a���?�?�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?      �?        333333�?�������?              �?/�袋.�?F]t�E�?              �?�������?�������?      �?                      �?w�qG��?⎸#��?              �?�������?333333�?      �?        �m۶m��?%I�$I��?              �?]t�E�?t�E]t�?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?      �?                      �?              �?UUUUUU�?�������?]t�E]�?�E]t��?֔5eMY�?�5eMYS�?�i��F�?	�=����?              �?I�$I�$�?۶m۶m�?�������?333333�?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?�q�q�?9��8���?      �?      �?              �?      �?              �?              �?        ى�؉��?�N��N��?              �?��y��y�?�a�a�?      �?      �?              �?      �?      �?      �?      �?      �?                      �?              �?�������?�������?      �?                      �?R���Q�?���Q��?F�:�$�?��KWm�?�S�<%��?pX���o�?,Q��+�?jW�v%j�?۶m۶m�?�$I�$I�?              �?      �?      �?�������?UUUUUU�?              �?      �?        �������?333333�?      �?      �?      �?                      �?      �?      �?              �?      �?        �������?�������?(�����?�5��P�?�$I�$I�?n۶m۶�?              �?      �?      �?      �?                      �?              �?      �?        �7��Mo�?d!Y�B�?�������?�������?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        �؉�؉�?;�;��?      �?        <<<<<<�?�?              �?      �?      �?�������?�?      �?        5�rO#,�?�{a���?]t�E]�?F]t�E�?              �?ffffff�?333333�?ZZZZZZ�?�������?      �?        ى�؉��?�؉�؉�?]t�E�?F]t�E�?              �?      �?                      �?              �?      �?        ��h����?��\���?      �?        ��S	�?��1����?      �?      �?�������?�������?l(�����?(������?۶m۶m�?�$I�$I�?�������?�������?�q�q�?9��8���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?              �?      �?              �?                      �?[k���Z�?�RJ)���?��(��(�?�\�\�?�����F�?W�+�ɵ?�������?�?      �?        ]t�E]�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        r�q��?9��8���?�c�1��?�s�9��?b'vb'v�?;�;��?�E]t��?]t�E]�?      �?      �?333333�?ffffff�?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?9��8���?�q�q�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?	�%����?h/�����?      �?              �?      �?              �?      �?              �?              �?        ��O ���?��`����?GS��r�?�b��7�?�������?�������?333333�?ffffff�?      �?      �?              �?      �?                      �?      �?        �o�z2~�?�@�6�?>���>�?|���?              �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?              �?              �?      �?              �?      �?        333333�?333333�?      �?      �?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        �5��P�?(�����?�k(���?(�����?n۶m۶�?�$I�$I�?�������?�������?      �?                      �?      �?        �������?�������?      �?      �?              �?      �?              �?              �?              �?      �?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJP�dhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM!hjh))��}�(h,h/h0M!��h2h3h4hph<�h=Kub������       X                    �?ʡ�;S��?�           8�@               S                    @�z�G��?�            @o@              :                   @B@��Q���?�             n@                                  �?
��^���?r            @g@                                ��.@     ��?)             P@                                  P,@�4�����?             ?@                                  �?�J�4�?             9@        ������������������������       �                     @        	       
                 ���@z�G�z�?             4@        ������������������������       �                      @                                �|�9@�����H�?             2@        ������������������������       �                     @                                   �?8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �@@               9                   �?@�̚��?I            �^@              2                 м�9@���|���?>            �X@                                  @�w��#��?"             I@        ������������������������       �                     @                                P�@p�v>��?            �G@                                   �?      �?              @                                 �7@����X�?             @        ������������������������       �                     @                                �&B@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?               '                     @x�����?            �C@                                    5@      �?              @        ������������������������       �                      @        !       &                   �<@�q�q�?             @       "       #                   �'@���Q��?             @        ������������������������       �                      @        $       %                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        (       )                   �9@`Jj��?             ?@       ������������������������       �        
             5@        *       1                    �?z�G�z�?             $@       +       ,                 @3�@���Q��?             @        ������������������������       �                     �?        -       0                 �|Y>@      �?             @       .       /                 pf&(@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        3       8                     @��<D�m�?            �H@       4       5                    �?`Ql�R�?            �G@       ������������������������       �                    �A@        6       7                    @�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     7@        ;       R                 �D�H@��}*_��?!             K@       <       I                   �G@և���X�?            �A@       =       B                    �? �o_��?             9@        >       A                   @F@�eP*L��?             &@       ?       @                   �,@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        C       D                 ��T?@@4և���?             ,@       ������������������������       �                     "@        E       F                    �?z�G�z�?             @        ������������������������       �                      @        G       H                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        J       O                     �?z�G�z�?             $@       K       L                   �H@r�q��?             @        ������������������������       �                     @        M       N                    K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        P       Q                   �*@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        T       U                 ��T?@ףp=
�?             $@        ������������������������       �                     @        V       W                    %@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        Y       �                 ��i=@�.����?           �|@       Z       _                    @`}C=|�?�            �u@        [       ^                    @r�q��?             @        \       ]                 �(\�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        `       �                   �4@��(�?�            0u@        a       d                     @�rF���?&            �K@        b       c                    &@      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        e       h                    �?��|�5��?             �G@        f       g                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        i       ~                    �?r�q��?             E@       j       {                    �?8�Z$���?            �C@       k       x                    �?��hJ,�?             A@       l       w                   �2@��a�n`�?             ?@        m       t                   �1@�z�G��?	             $@       n       s                   �0@؇���X�?             @        o       p                 pf�@�q�q�?             @        ������������������������       �                     �?        q       r                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        u       v                 ��Y @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        y       z                  s�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        |       }                 032@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @               �                    #@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�7�2�?�            �q@       �       �                   �F@����?�            �p@       �       �                    �?�s�c���?�            �l@        �       �                     @��a�n`�?             ?@        ������������������������       �                     @        �       �                 �|Y=@R�}e�.�?             :@        �       �                   �6@�q�q�?             "@        ������������������������       �                     �?        �       �                 �0@      �?              @       �       �                    �?      �?             @       �       �                   @:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   @@�IєX�?             1@       �       �                 �|�=@�C��2(�?             &@       �       �                 ���@؇���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��$:@DGr���?�             i@       �       �                     �?����W�?|            `h@        ������������������������       �                     @        �       �                 ���@�:nR&y�?x            �g@        ������������������������       �                     5@        �       �                 ���@0u��Fs�?k             e@        ������������������������       �                      @        �       �                   �<@�8��?j            �d@        ������������������������       �        "            �K@        �       �                   @@@ �Cc}�?H             \@       �       �                    �?      �?3             T@       �       �                 ��@���!���?2            �S@        ������������������������       �                     4@        �       �                    �?@�r-��?'            �M@        ������������������������       �                     @        �       �                    �?�2����?$            �K@       �       �                 �|�=@�iʫ{�?#            �J@       �       �                 ��) @tk~X��?             B@       �       �                  sW@�8��8��?             8@        ������������������������       �      �?             @        ������������������������       �                     4@        �       �                     @�q�q�?             (@        �       �                 �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    (@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �@�t����?             1@        �       �                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�@��S�ۿ?             .@        �       �                 �?�@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     �?        �       �                     @      �?             @@        �       �                   �3@��S�ۿ?
             .@       �       �                 `fF)@�����H�?             "@        ������������������������       �                     �?        �       �                   @D@      �?              @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                   �B@�IєX�?             1@        ������������������������       �                     @        �       �                 @3�@ףp=
�?             $@        �       �                   �C@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 X�,@@���Q��?             @        ������������������������       �                     �?        �       �                 03k:@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     D@        �       �                    �?�θ�?
             *@        ������������������������       �                     �?        �       �                 �|Y?@      �?	             (@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �                          �R@Ц����?@             ]@       �                          @d}h��??             \@       �                          E@X&$�E�?6            �X@       �                          �?     ��?#             P@       �       �                     @�q�����?             I@       �       �                    �?~�4_�g�?             F@        �       �                  Y>@�z�G��?
             4@        ������������������������       �                     @        �       �                 �|Y<@      �?             0@        ������������������������       �                     @        �       �                 X�,@@���Q��?             $@        ������������������������       �                     @        �       �                   �A@�q�q�?             @        ������������������������       �                      @        �       �                 @�Cq@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @A@�q�q�?             8@       �       �                    �?�㙢�c�?             7@       �       �                 �|Y>@      �?
             0@       �       �                     �?����X�?	             ,@       �       �                   �;@�	j*D�?             *@        ������������������������       �                     �?        �       �                 �|�<@      �?             (@        �       �                 `f�D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �>@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �                           >@r�q��?             @       �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @              	                   �?����X�?             ,@                                 �?"pc�
�?             &@                               �4@z�G�z�?             $@        ������������������������       �                     @                              �̾w@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        
                         �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 �?(N:!���?            �A@        ������������������������       �        	             3@                              0��M@      �?
             0@                                �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?8�Z$���?             *@                               �G@�q�q�?             @        ������������������������       �                     @                                 �?�q�q�?             @                             @��V@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                              ���A@$�q-�?	             *@                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M!KK��h2h3h4hVh<�h=Kub������������N���I5�?d�~`l��?333333�?ffffff�?�������?333333�?��~���?X`��?      �?      �?��RJ)��?���Zk��?{�G�z�?�z�G��?              �?�������?�������?      �?        �q�q�?�q�q�?              �?;�;��?;�;��?              �?      �?              �?                      �?�u�y���??�%C���?F]t�E�?]t�E]�?��Q��?��(\���?              �?ڨ�l�w�?L� &W�?      �?      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?��o��o�?�A�A�?      �?      �?              �?UUUUUU�?UUUUUU�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?���{��?�B!��?      �?        �������?�������?333333�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        և���X�?��S�r
�?W�+�ɕ?}g���Q�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?B{	�%��?_B{	�%�?�$I�$I�?۶m۶m�?
ףp=
�?�Q����?]t�E�?t�E]t�?      �?      �?      �?                      �?      �?        n۶m۶�?�$I�$I�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?              �?�������?�������?      �?        �������?�������?              �?      �?        �/R��?�@���'�?��"9��?�tS�?UUUUUU�?�������?      �?      �?              �?      �?                      �?�Ź�Q�?�8�1�s�?yJ���?�־a��?      �?      �?      �?      �?      �?        br1���?x6�;��?�������?�������?              �?      �?        �������?UUUUUU�?;�;��?;�;��?KKKKKK�?�������?�s�9��?�c�1Ƹ?ffffff�?333333�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ����.��?�
��V�?�]�\�*�?�e�?�����?�cj`?�c�1��?�s�9��?      �?        'vb'vb�?�;�;�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?                      �?�?�?]t�E�?F]t�E�?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?              �?        H�z�G�?��(\�µ?>۳=۳�?&a&a�?      �?        Fڱa��?�-q��ܲ?      �?         s�n_Y�?g\�5�?              �?y�oqZ��?7Āt,e�?      �?        %I�$I��?۶m۶m�?      �?      �?��	�Z�?T:�g *�?      �?        'u_�?��c+���?      �?        ��7�}��?� O	��?
�[���?�琚`��?r�q��?9��8���?UUUUUU�?UUUUUU�?      �?      �?      �?        �������?�������?      �?      �?      �?                      �?      �?      �?              �?      �?        <<<<<<�?�?      �?      �?      �?                      �?�������?�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?                      �?      �?      �?�������?�?�q�q�?�q�q�?      �?              �?      �?      �?              �?      �?      �?        �?�?      �?        �������?�������?      �?      �?UUUUUU�?UUUUUU�?      �?              �?        �������?333333�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?        ى�؉��?�؉�؉�?      �?              �?      �?      �?      �?              �?      �?              �?        �4�rO#�?�{a��?�m۶m��?�$I�$I�?b�ΐ���?;Cb�ΐ�?      �?      �?�p=
ף�?���Q��?/�袋.�?��.���?333333�?ffffff�?              �?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?UUUUUU�?�������?�7��Mo�?d!Y�B�?      �?      �?�m۶m��?�$I�$I�?vb'vb'�?;�;��?              �?      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?              �?              �?              �?                      �?UUUUUU�?�������?      �?      �?              �?      �?                      �?�$I�$I�?�m۶m��?F]t�E�?/�袋.�?�������?�������?              �?�������?333333�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        |�W|�W�?�A�A�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?        �؉�؉�?;�;��?      �?      �?              �?      �?              �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�g?BhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       Z                    �?S*f���?�           8�@               ?                 �|�=@�-�����?�             n@                                   @NU��b��?`            �a@                                   �?      �?'             P@                                  �?P���Q�?             D@        ������������������������       �        
             ,@                                   9@$�q-�?             :@                                 �3@8�Z$���?             *@        	       
                   �'@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     *@        ������������������������       �                     8@                                    �?rOP\6�?9            @S@                                   �?      �?             @@                               ���@���7�?             6@                                �|Y5@�q�q�?             @        ������������������������       �                     �?                                �Y�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@                                `�@1@�z�G��?             $@                                   �?      �?             @                                  �?�q�q�?             @        ������������������������       �                     �?                                �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        !       :                    �?X�<ݚ�?!            �F@       "       #                    &@4���C�?            �@@        ������������������������       �                     @        $       5                   �;@      �?             <@       %       &                 P��@j���� �?             1@        ������������������������       �                     @        '       0                   �9@      �?             ,@       (       )                 @33"@      �?              @        ������������������������       �                     @        *       /                   �6@���Q��?             @       +       ,                 ��,#@      �?             @        ������������������������       �                     �?        -       .                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        1       4                   �:@�q�q�?             @       2       3                 pf(@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        6       9                    �?���|���?             &@       7       8                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ;       <                    �?�8��8��?	             (@        ������������������������       �                     @        =       >                    @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        @       S                     @�ڊ�e��?>             Y@       A       D                 ���&@�ƫ�%�?6            @V@        B       C                   �J@      �?             @       ������������������������       �                     @        ������������������������       �                     @        E       F                   �B@ Df@��?3            �T@        ������������������������       �                     A@        G       H                     �?@9G��?             �H@       ������������������������       �                     ?@        I       N                    �?�����H�?	             2@        J       M                   �*@      �?              @        K       L                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        O       R                    �?ףp=
�?             $@        P       Q                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        T       Y                   @C@���|���?             &@       U       V                    �?      �?              @        ������������������������       �                     �?        W       X                   �>@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        [       �                 `�X.@Έx�Ȝ�?.           `}@       \       q                 �?�@���o[�?�            �q@        ]       p                    �?г�wY;�?\             a@       ^       c                   �6@ ����O�?Y            ``@        _       `                   �5@�KM�]�?             3@       ������������������������       �                     .@        a       b                 03�@      �?             @        ������������������������       �                      @        ������������������������       �                      @        d       e                  ��@�h����?K             \@        ������������������������       �        %            �J@        f       o                 �?$@���#�İ?&            �M@        g       j                 ��@�C��2(�?             6@       h       i                 �|Y=@�IєX�?
             1@        ������������������������       �                     �?        ������������������������       �        	             0@        k       l                 �|�;@z�G�z�?             @        ������������������������       �                     @        m       n                 �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �B@        ������������������������       �                     @        r       �                    �?�npº��?_            �b@       s       �                    �?���H��?T            �`@       t       �                     @ףp=
�?R            @`@        u       x                    5@���7�?             F@        v       w                    &@r�q��?             @       ������������������������       �      �?              @        ������������������������       �                     @        y       �                   @A@P�Lt�<�?             C@       z       {                 `fF)@�}�+r��?             3@        ������������������������       �                     @        |                        ��,@�8��8��?	             (@       }       ~                    @@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        �       �                    �?���tT��?4            �U@        ������������������������       �                     �?        �       �                 �|Y=@|�M���?3            @U@        �       �                   �:@�������?             F@       �       �                 0S5 @$G$n��?            �B@        �       �                   �3@     ��?             0@        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     5@        �       �                   �;@և���X�?             @        ������������������������       �                     @        �       �                   �<@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @C@������?            �D@       �       �                 ��) @      �?             @@       ������������������������       �                     5@        �       �                 ��y @�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 @3�@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �4@�E��ӭ�?             2@        ������������������������       �                     @        ������������������������       �                     *@        �       �                    #@:v�S��?s            �f@        �       �                    @$��m��?             :@       ������������������������       �        	             .@        �       �                    @"pc�
�?             &@       �       �                    @�q�q�?             @       �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                 ���A@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?������?b            �c@        �       �                    I@      �?!             E@       �       �                 �̾w@��
ц��?            �C@       �       �                    �?��
P��?            �A@       �       �                    �?b�2�tk�?             2@       �       �                 `f�A@�eP*L��?
             &@       �       �                      @����X�?             @       �       �                 X�,@@z�G�z�?             @       �       �                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �7@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    3@j���� �?             1@        ������������������������       �                     �?        �       �                    �?      �?             0@        �       �                     �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y>@և���X�?             @       �       �                     @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `ff:@�㙢�c�?A            �\@        ������������������������       �                     ?@        �       �                 03�>@���N8�?-             U@        �       �                    K@��>4և�?             <@       �       �                    �?�\��N��?             3@       �       �                   @>@����X�?             ,@       �       �                   �<@X�<ݚ�?             "@        ������������������������       �                      @        �       �                 `f�;@և���X�?             @       �       �                 X��B@      �?             @        ������������������������       �                     �?        �       �                   @G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        �       �                   @=@�q�q�?             @        ������������������������       �                     �?        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �Q@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                    J@�X�C�?             L@       �       �                    �?�������?             F@       �       �                 03�U@     ��?             @@       �       �                     @V�a�� �?             =@       �       �                 03�I@�㙢�c�?             7@        ������������������������       �                      @        �       �                 `�iJ@������?             .@        ������������������������       �                      @        �       �                   @K@8�Z$���?             *@        �       �                    7@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    ;@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     (@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������H�7�?=�o�a��?�>�>�?�T��T��?qJ��O$�?d-C���?      �?      �?�������?ffffff�?              �?;�;��?�؉�؉�?;�;��?;�;��?      �?      �?              �?      �?                      �?              �?              �?dj`��?��O����?      �?      �?F]t�E�?�.�袋�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?333333�?ffffff�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?r�q��?�q�q�?'�l��&�?m��&�l�?              �?      �?      �?ZZZZZZ�?�������?              �?      �?      �?      �?      �?      �?        �������?333333�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?�������?333333�?              �?      �?                      �?]t�E]�?F]t�E�?۶m۶m�?�$I�$I�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?              �?      �?        
ףp=
�?��Q��?�as�ì?��x�3�?      �?      �?              �?      �?        ��k���?c��7�:�?              �?9/���?������?              �?�q�q�?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?      �?              �?      �?                      �?F]t�E�?]t�E]�?      �?      �?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?        �t�SY�?�-z���?�oAi6�?���L�?�?�?����?qBJ�eD�?�k(���?(�����?      �?              �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?        ��N��?'u_[�?]t�E�?F]t�E�?�?�?              �?      �?        �������?�������?      �?              �?      �?              �?      �?              �?              �?        �2n���?�4G�#��?h	&�?���̾?�������?�������?�.�袋�?F]t�E�?�������?UUUUUU�?      �?      �?      �?        ���k(�?(�����?�5��P�?(�����?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?              �?        ����/��?�}A_�?      �?        �������?�������?t�E]t�?/�袋.�?к����?���L�?      �?      �?              �?      �?              �?        ۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?p>�cp�?������?      �?      �?      �?        ]t�E�?F]t�E�?              �?      �?        �q�q�?�q�q�?              �?      �?                      �?�q�q�?r�q��?              �?      �?        '<�ߠ��?��Y@�H�?vb'vb'�?�N��N��?              �?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?333333�?�������?      �?              �?      �?              �?      �?              �?              �?        �����?X�˟��?      �?      �?�؉�؉�?�;�;�?PuPu�?_�_��?�8��8��?9��8���?t�E]t�?]t�E�?�$I�$I�?�m۶m��?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?      �?        �m۶m��?�$I�$I�?              �?      �?        ZZZZZZ�?�������?      �?              �?      �?�q�q�?9��8���?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?                      �?      �?        �7��Mo�?d!Y�B�?      �?        �a�a�?��y��y�?۶m۶m�?I�$I�$�?�5��P�?y�5���?�$I�$I�?�m۶m��?�q�q�?r�q��?              �?�$I�$I�?۶m۶m�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?      �?        �q�q�?�q�q�?      �?                      �?�m۶m��?%I�$I��?t�E]t�?/�袋.�?      �?      �?��{a�?a���{�?�7��Mo�?d!Y�B�?      �?        wwwwww�?�?              �?;�;��?;�;��?333333�?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ1�.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM-hjh))��}�(h,h/h0M-��h2h3h4hph<�h=Kub������                        x#J@� ��4d�?�           8�@              ]                    �?�~���?|           Ђ@               @                    �?�y��<��?`            `c@                                   �?4uj�w��?D            @\@                                ��";@��<b���?             7@        ������������������������       �                     �?                                ��4=@"pc�
�?             6@        ������������������������       �                     @        	                          �@@������?
             .@        
                        �|�=@      �?             @                               03SA@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                 �>@�C��2(�?             &@        ������������������������       �                     @                                p�i@@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?���Q��?6            �V@                                ��*@�<ݚ�?             ;@                               �|Y8@���}<S�?             7@        ������������������������       �                     "@                                    @؇���X�?
             ,@        ������������������������       �                      @                                 ��@r�q��?             (@                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                1                 �|Y=@���N8�?$            �O@        !       "                     @j���� �?
             1@        ������������������������       �                      @        #       $                 ���@�q�q�?	             .@        ������������������������       �                      @        %       0                    �?�θ�?             *@       &       )                   @@r�q��?             (@        '       (                   �5@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        *       /                    �?؇���X�?             @       +       ,                 ��*@r�q��?             @        ������������������������       �                     �?        -       .                   �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        2       9                    �?�q��/��?             G@       3       8                   @@�����?             5@       4       7                 �|�=@r�q��?	             (@       5       6                 ���@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     "@        :       ;                 ���@H%u��?             9@        ������������������������       �                     @        <       ?                 X��A@r�q��?
             2@       =       >                   @'@@�0�!��?	             1@       ������������������������       �z�G�z�?             .@        ������������������������       �                      @        ������������������������       �                     �?        A       V                 `v�9@�G��l��?             E@       B       I                    �?J�8���?             =@       C       H                 ��.@������?
             .@        D       E                   �-@�q�q�?             @        ������������������������       �                     @        F       G                 �|Y6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        J       S                    �?և���X�?	             ,@       K       L                     @X�<ݚ�?             "@        ������������������������       �                     �?        M       P                    �?      �?              @       N       O                 �&�)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Q       R                   `3@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        T       U                   �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        W       X                     �?�θ�?	             *@        ������������������������       �                     �?        Y       Z                  �=@r�q��?             (@        ������������������������       �                     @        [       \                   �3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ^       �                    �?节>t�?           �{@        _       �                    �?��rf�B�?O            @_@       `       �                    @�
I���?D             [@       a       t                 `f�$@�O��i�?@            �Y@        b       o                    �?f���M�?             ?@       c       j                    7@�û��|�?             7@       d       i                   �4@�q�q�?             (@       e       h                 @3"@և���X�?             @       f       g                 P��@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        k       l                 �|Y>@�C��2(�?             &@        ������������������������       �                     @        m       n                    A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        p       s                    �?      �?              @       q       r                    4@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        u       �                   �K@r�q��?.             R@       v                            @�~t��?,            @Q@       w       ~                    6@      �?             H@        x       }                   �;@��2(&�?             6@        y       z                   �'@և���X�?             @        ������������������������       �                     @        {       |                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             .@        ������������������������       �                     :@        �       �                    @�q�q�?             5@        ������������������������       �                      @        �       �                 �|�<@��
ц��?	             *@        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                    �?����X�?             @       �       �                    �?r�q��?             @       �       �                 �|Y>@�q�q�?             @        ������������������������       �                     �?        �       �                 03�1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���3@�IєX�?             1@        �       �                   `2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             .@        �       �                    �?Ї	{�k�?�             t@       �       �                   @R@ףp=
�?�             r@       �       �                 ��$:@A��Tf�?�            r@       �       �                    �?����?�            `o@       �       �                 �?�@��Au5a�?�            �k@        �       �                 �?$@X;��?8            @V@       �       �                     @0G���ջ?"             J@        ������������������������       �                     @        �       �                 �|Y>@���.�6�?             G@       �       �                 ���@     ��?             @@       �       �                 ���@ �q�q�?             8@        �       �                    7@ףp=
�?             $@        ������������������������       �                     @        �       �                   �8@r�q��?             @        �       �                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             ,@        �       �                 �|�;@      �?              @        ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �        	             ,@        ������������������������       �                    �B@        �       �                   �@@�8��8��?R            �`@       �       �                   �2@h�a��?;            @X@        �       �                   �1@8�Z$���?
             *@       �       �                 pf� @ףp=
�?             $@        ������������������������       �      �?              @        ������������������������       �                      @        �       �                     @�q�q�?             @        ������������������������       �                     �?        �       �                 ��Y @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�!@h�����?1             U@        �       �                 ��) @��p\�?            �D@       ������������������������       �                     ;@        �       �                    8@d}h���?             ,@        ������������������������       �                     @        �       �                 �|�>@      �?              @       �       �                 �|Y<@      �?             @        ������������������������       �                      @        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �E@        �       �                     @b�h�d.�?            �A@       �       �                   �*@�<ݚ�?             2@       �       �                    G@���Q��?             $@        �       �                   �'@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @D@�t����?
             1@        �       �                 @3�@      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     >@        �       �                     �?p�ݯ��?             C@       �       �                 �|Y>@؀�:M�?            �B@        �       �                   `@@      �?             (@       �       �                 `fF<@ףp=
�?             $@        �       �                 �|�<@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    @@z�G�z�?             9@       �       �                 03k:@�q�q�?             .@        ������������������������       �                     �?        �       �                   �=@����X�?
             ,@       �       �                 `f�;@�θ�?	             *@       �       �                   �J@�q�q�?             "@        �       �                   @G@      �?             @        �       �                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    :@     ��?             @@       �       �                 ���'@X�Cc�?             ,@        ������������������������       �                     @        �       �                    )@      �?
             $@       �       �                 @3�4@r�q��?             @       ������������������������       �                     @        �       �                 ���7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�����H�?
             2@        �       �                    @�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 ��T?@؇���X�?             @       ������������������������       �                     @                                  @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @              $                    �? ��?�?F            @[@                                �?�+I�9��?<            @V@                                �?�g�y��?+             O@       ������������������������       �        %             K@                                 �?      �?              @        ������������������������       �                     �?        	                      Ъ�c@����X�?             @        
                         3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?l��
I��?             ;@                                �?�q�q�?             2@                                 �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @                                 �?X�<ݚ�?             "@                             `f�N@և���X�?             @                             ��9L@���Q��?             @                                7@      �?             @        ������������������������       �                     �?                                @K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @              #                  �G@�<ݚ�?             "@                                 �?      �?              @        ������������������������       �                     @        !      "                �̰f@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        %      ,                   �?z�G�z�?
             4@        &      +                  PQ@���Q��?             $@       '      (                   ;@X�<ݚ�?             "@        ������������������������       �                     @        )      *                   �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �*       h�h))��}�(h,h/h0M-KK��h2h3h4hVh<�h=Kub��������������`uv��?,J>��?�� [	��?�L�I�-�?���/Y��?�4�M�?�:Fq�c�?2�s�8�?��,d!�?��Moz��?              �?/�袋.�?F]t�E�?      �?        wwwwww�?�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?]t�E�?F]t�E�?      �?        �������?�������?              �?      �?        333333�?�������?�q�q�?9��8���?d!Y�B�?ӛ���7�?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?        �a�a�?��y��y�?ZZZZZZ�?�������?      �?        UUUUUU�?UUUUUU�?      �?        �؉�؉�?ى�؉��?UUUUUU�?�������?�������?�������?              �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?�������?              �?�������?�������?      �?                      �?              �?      �?        �B����?��Mozӻ?=��<���?�a�a�?�������?UUUUUU�?9��8���?�q�q�?      �?        333333�?�������?      �?              �?        )\���(�?���Q��?      �?        �������?UUUUUU�?ZZZZZZ�?�������?�������?�������?      �?              �?        ��y��y�?1�0��?|a���?�rO#,��?�?wwwwww�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?۶m۶m�?�$I�$I�?r�q��?�q�q�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?      �?                      �?�������?�������?      �?                      �?ى�؉��?�؉�؉�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �����D�?�y����?�A`��"�?;�O��n�?�^B{	��?��^B{	�?��,��?�����?��RJ)��?��Zk���?8��Moz�?��,d!�?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?              �?]t�E�?F]t�E�?      �?              �?      �?              �?      �?              �?      �?�m۶m��?�$I�$I�?              �?      �?              �?        UUUUUU�?�������?)�3J���?�s��\�?      �?      �?t�E]t�?��.���?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?�;�;�?�؉�؉�?      �?              �?      �?              �?�$I�$I�?�m۶m��?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �?�?      �?      �?      �?                      �?      �?        6�l�?�O���?�������?�������?��"�O��?U��6�͸?Pv�`7�?���Ɏ�?�����?�7�7�?�u�{���?�E(B�?vb'vb'�?�؉�؉�?      �?        ���7���?Y�B��?      �?      �?�������?UUUUUU�?�������?�������?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?              �?              �?      �?      �?        333333�?�������?      �?              �?        UUUUUU�?UUUUUU�?�D�a�Y�?���Id�?;�;��?;�;��?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �m۶m��?�$I�$I�?�]�ڕ��?��+Q��?      �?        I�$I�$�?۶m۶m�?      �?              �?      �?      �?      �?              �?      �?      �?              �?      �?              �?              �?        ;��:���?_�_��?9��8���?�q�q�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        <<<<<<�?�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?              �?        ^Cy�5�?Cy�5��?E>�S��?v�)�Y7�?      �?      �?�������?�������?      �?      �?              �?      �?                      �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?�m۶m��?�$I�$I�?ى�؉��?�؉�؉�?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?                      �?      �?              �?                      �?      �?              �?                      �?      �?      �?%I�$I��?�m۶m��?      �?              �?      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        �q�q�?�q�q�?]t�E�?F]t�E�?              �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���]8��?߅���]�?�as�ü?�3��g�?�B!��?��{���?              �?      �?      �?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?h/�����?Lh/����?UUUUUU�?UUUUUU�?�q�q�?9��8���?      �?                      �?�q�q�?r�q��?�$I�$I�?۶m۶m�?�������?333333�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�q�q�?9��8���?      �?      �?              �?�������?�������?              �?      �?              �?        �������?�������?333333�?�������?r�q��?�q�q�?              �?�������?UUUUUU�?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg�)hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM!hjh))��}�(h,h/h0M!��h2h3h4hph<�h=Kub������       �                  x#J@���?Y��?�           8�@                                  @���>�?}           ��@                                   @$G$n��?            �B@                                  @�<ݚ�?             2@       ������������������������       �        
             ,@        ������������������������       �                     @                                   @�}�+r��?             3@       ������������������������       �                     .@        	       
                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?               a                    �?d[��8X�?g           x�@               R                    �?���(�_�?o            �e@              !                     @�%o��?V            �`@                                  �B@�C��2(�?&            �K@                                  6@P�Lt�<�?             C@                                   �?      �?             0@       ������������������������       �        	             ,@                                ��m1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@                                 03{;@������?             1@                                 �C@     ��?
             0@        ������������������������       �                      @                                    �?@4և���?	             ,@        ������������������������       �                     @                                  @F@�C��2(�?             &@                                  �E@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        "       I                    �?V�K/��?0            �S@       #       8                    �?�xGZ���?(            �Q@       $       )                    �?��J�fj�?            �B@        %       (                 �&�@�r����?             .@        &       '                 0��@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        *       /                   �7@���|���?             6@        +       ,                   �3@      �?              @        ������������������������       �                     �?        -       .                 ��|!@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        0       7                   &@d}h���?             ,@       1       6                   �@�8��8��?             (@        2       3                   �9@z�G�z�?             @        ������������������������       �                     @        4       5                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        9       B                    �?�'�=z��?            �@@        :       =                   �-@X�Cc�?             ,@        ;       <                   �,@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        >       ?                 �|Y6@�����H�?             "@        ������������������������       �                      @        @       A                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        C       F                 �|�;@D�n�3�?             3@        D       E                 P�@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        G       H                 03�1@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        J       M                    �?X�<ݚ�?             "@        K       L                 ��*@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        N       Q                 �A7@�q�q�?             @       O       P                 ���1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        S       T                     @�99lMt�?            �C@        ������������������������       �                     "@        U       \                  Y3@r�q��?             >@        V       [                    �?�q�q�?             @       W       X                 ���&@�q�q�?             @        ������������������������       �                     �?        Y       Z                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ]       ^                    @ �q�q�?             8@       ������������������������       �        
             1@        _       `                   @C@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        b       }                     �?�ը
q��?�             x@        c       v                  �>@6�iL�?"            �M@       d       u                    �?�eP*L��?            �@@       e       l                    �?�g�y��?             ?@        f       k                   @G@����X�?             @       g       j                 �ܵ<@r�q��?             @        h       i                 ��";@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        m       t                   @>@�q�q�?             8@       n       o                   �<@@�0�!��?	             1@        ������������������������       �                      @        p       q                 03:@��S�ۿ?             .@        ������������������������       �                     "@        r       s                 03k:@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        w       |                    �? ��WV�?             :@       x       {                 �|�<@�nkK�?             7@        y       z                 `f�D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        ������������������������       �                     @        ~       �                     @H�` |�?�            pt@               �                    4@ ��Ou��?3            �S@        �       �                    &@�<ݚ�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                 �|Y=@�nkK�?.            @Q@        ������������������������       �                     3@        �       �                    �? "��u�?"             I@       �       �                    �?���.�6�?             G@        ������������������������       �                     @        �       �                    �?��(\���?             D@       �       �                 `f�)@�#-���?            �A@        ������������������������       �        	             .@        �       �                   �*@R���Q�?             4@       �       �                 �|�=@�z�G��?	             $@        ������������������������       �                     �?        �       �                    @@�<ݚ�?             "@        ������������������������       �                      @        �       �                   �A@����X�?             @        ������������������������       �                     �?        �       �                   @D@r�q��?             @        ������������������������       �                      @        �       �                    G@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     @        �       �                   @@@H�@>��?�             o@       �       �                    �?"����U�?�            @i@        �       �                    �?��N`.�?&            �K@       �       �                    �?z�G�z�?             D@       �       �                   �+@�+e�X�?             9@       �       �                 �|Y=@�q�q�?             8@        �       �                 ��y@      �?              @        ������������������������       �                      @        �       �                   @9@�q�q�?             @        ������������������������       �                     @        �       �                   @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|�=@      �?             0@       �       �                 ���@�8��8��?	             (@        ������������������������       �                     @        �       �                   @@      �?              @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                  ��@�r����?             .@        ������������������������       �                      @        ������������������������       �����X�?             @        �       �                    �?�q�q�?
             .@       �       �                 03�-@�<ݚ�?             "@        �       �                    3@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 03�7@      �?             @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �>@\�JЂ.�?a            `b@       �       �                    #@���	���?\             a@        �       �                     @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?���D�k�?Y            �`@       �       �                 @3�@L�'�7��?L            @]@       �       �                   �7@P�2E��?-            @P@        ������������������������       �                     9@        �       �                   �8@��(\���?             D@        �       �                 `fF@����X�?             @        �       �                 �&b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|�<@Pa�	�?            �@@        ������������������������       �                     "@        �       �                 �|�=@ �q�q�?             8@       �       �                  sW@�nkK�?             7@        �       �                 pf�@�C��2(�?             &@       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     (@        ������������������������       �                     �?        �       �                   �2@8�Z$���?             J@        �       �                 ��Y @      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                 0S%"@�Ra����?             F@       �       �                 ��) @�GN�z�?             6@       �       �                   �5@��S�ۿ?             .@        ������������������������       �      �?              @        ������������������������       �        	             *@        �       �                    8@և���X�?             @        ������������������������       �                      @        �       �                 �|Y<@z�G�z�?             @        ������������������������       �                     �?        �       �                 pf� @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             6@        ������������������������       �                     0@        �       �                   �?@���Q��?             $@        ������������������������       �                      @        �       �                   �@      �?              @        ������������������������       �                     �?        �       �                 �?�@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                    �G@        �                           @�㙢�c�?F            �\@       �                          �?r�q��?E            �\@        �       �                    �?ȵHPS!�?             J@       �       �                      @h�����?             <@       ������������������������       �                     8@        �       �                    >@      �?             @       �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �                           �?�q�q�?             8@        �       �                    �?z�G�z�?             $@        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                �B@d}h���?             ,@       ������������������������       �                     $@                                 �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                 �?�z�6�?&             O@              
                  �2@      �?             @@              	                ��e@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @                              �UcV@8�Z$���?             :@        ������������������������       �                     ,@                                 E@�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @                                 �?r�q��?             >@                                T@PN��T'�?             ;@                               �M@      �?             0@                                �?z�G�z�?             .@       ������������������������       �                     "@                                 A@      �?             @                             `f�K@      �?             @                                7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0M!KK��h2h3h4hVh<�h=Kub��������������� 3��?@Bx���?xR��y��?[���?���L�?к����?�q�q�?9��8���?              �?      �?        (�����?�5��P�?              �?      �?      �?              �?      �?        �w����?��"��?�wK�?��?DZ/`��?\�՘H�?���[��?F]t�E�?]t�E�?(�����?���k(�?      �?      �?              �?      �?      �?              �?      �?                      �?�?xxxxxx�?      �?      �?      �?        �$I�$I�?n۶m۶�?              �?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �Z܄��?�ґ=�?�A�A�?�_�_�?к����?�"�u�)�?�?�������?      �?      �?              �?      �?                      �?]t�E]�?F]t�E�?      �?      �?      �?        �$I�$I�?�m۶m��?              �?      �?        I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?              �?                      �?|���?|��|�?�m۶m��?%I�$I��?�������?�������?              �?      �?        �q�q�?�q�q�?              �?�$I�$I�?۶m۶m�?      �?                      �?l(�����?(������?]t�E�?F]t�E�?              �?      �?              �?      �?              �?      �?        r�q��?�q�q�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        5H�4H��?�o��o��?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�������?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        ��
��[�?����?ylE�pR�?'u_[�?t�E]t�?]t�E�?�B!��?��{���?�$I�$I�?�m۶m��?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?�������?ZZZZZZ�?�������?              �?�������?�?      �?        �������?UUUUUU�?              �?      �?                      �?      �?        O��N���?;�;��?�Mozӛ�?d!Y�B�?      �?      �?              �?      �?              �?              �?        _�/���?
��֢P�?.��-���?�i�i�?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?        �Mozӛ�?d!Y�B�?      �?        �G�z�?���Q��?���7���?Y�B��?      �?        �������?333333�?�A�A�?_�_�?      �?        333333�?333333�?ffffff�?333333�?              �?9��8���?�q�q�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?              �?              �?              �?        @R0����?�>����?e�F�t�?j䮟-�?��oX���?� O	��?�������?�������?R���Q�?���Q��?UUUUUU�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?      �?              �?                      �?�������?�?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?�q�q�?9��8���?      �?      �?              �?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?        W�7�L�?gG-B���?V��,���?P�9��J�?      �?      �?              �?      �?        �՝VwZ�?�RKE,�?�������?���?_�^��?z�z��?      �?        �������?333333�?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        |���?|���?      �?        �������?UUUUUU�?�Mozӛ�?d!Y�B�?]t�E�?F]t�E�?      �?              �?      �?      �?              �?        ;�;��?;�;��?      �?      �?              �?      �?        ]t�E]�?]t�E�?�袋.��?]t�E�?�������?�?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?      �?              �?      �?              �?              �?        333333�?�������?              �?      �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?        d!Y�B�?�7��Mo�?UUUUUU�?�������?�؉�؉�?��N��N�?�$I�$I�?�m۶m��?              �?      �?      �?      �?      �?              �?      �?                      �?�������?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        ۶m۶m�?I�$I�$�?              �?      �?      �?              �?      �?        �Zk����?J)��RJ�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?h/�����?&���^B�?      �?      �?�������?�������?              �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�]_AhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       X                 @3�"@^����[�?�           8�@                                   �?���B���?�            @p@                                   @$��m��?             J@                                  �?ҳ�wY;�?            �I@                                   �?      �?             8@        ������������������������       �                     @                                ���@�S����?             3@        ������������������������       �                      @        	       
                    �?�IєX�?             1@       ������������������������       �        
             0@        ������������������������       �                     �?                                   ;@X�<ݚ�?             ;@                                  �?b�2�tk�?             2@                                 �3@�q�q�?	             .@                                P��@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                pf� @z�G�z�?             $@                               P�@�����H�?             "@       ������������������������       �                     @                                  �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                P�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                �?� @�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                7                   @4@$�q-�?�             j@        !       &                    �?�������?             >@        "       %                    �?���Q��?             @       #       $                 �{@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        '       4                    �?z�G�z�?             9@       (       3                   �2@��s����?             5@        )       0                   �1@���|���?             &@       *       /                   �0@      �?              @       +       ,                 pf�@�q�q�?             @        ������������������������       �                      @        -       .                 pFD!@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        1       2                 ��Y @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             $@        5       6                    3@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        8       E                   �8@�;Y�&��?n            @f@        9       :                   �5@�t����?             A@        ������������������������       �                     (@        ;       <                    �?"pc�
�?             6@        ������������������������       �                      @        =       D                    �?ףp=
�?             4@       >       ?                   �7@�KM�]�?             3@       ������������������������       �                     (@        @       C                 `fF@����X�?             @        A       B                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        F       O                   �>@@ݚ)�?Z             b@       G       H                    �?@uvI��?@            �X@        ������������������������       �                     C@        I       N                   �;@ �.�?Ƞ?)             N@        J       K                   �:@$�q-�?	             *@       ������������������������       �                     &@        L       M                 �� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �G@        P       Q                      @���}<S�?             G@        ������������������������       �                     �?        R       W                   @@@�:�^���?            �F@        S       T                   �?@      �?              @        ������������������������       �                     �?        U       V                 P�@և���X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                    �B@        Y       �                  x#J@������?           0|@       Z       �                    �?�ܨ`�?�            u@        [       f                    �?�E����?U             b@        \       a                 ��.@������?             >@        ]       `                 �|Y<@�eP*L��?             &@       ^       _                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        b       e                     �?�KM�]�?             3@        c       d                   �H@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@        g       �                    @�q�q�?C            �\@       h       �                    @F��L�?A            @[@       i       �                     @��wy���?7             W@       j                           :@ ,��-�?%            �M@       k       v                    �?�C��2(�?             F@       l       u                   �J@�FVQ&�?            �@@       m       t                   �*@      �?             @@       n       o                   �'@���N8�?             5@        ������������������������       �                     @        p       s                    �?      �?             0@       q       r                    B@@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        w       z                    6@"pc�
�?	             &@        x       y                   �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        {       ~                    �?�����H�?             "@       |       }                   �E@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             .@        �       �                    �?�eP*L��?            �@@        �       �                    '@j���� �?             1@        ������������������������       �                     @        �       �                   �@@�θ�?             *@       ������������������������       �                     "@        �       �                 `f�/@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?     ��?
             0@       �       �                   �;@���!pc�?             &@       ������������������������       �                     @        �       �                 `fv1@���Q��?             @        ������������������������       �                      @        �       �                 `fV6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    1@���Q��?             @       �       �                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?@�0�!��?
             1@        ������������������������       �                      @        �       �                 ��T?@��S�ۿ?	             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    '@�%����?|             h@        �       �                   �C@      �?             8@       �       �                    @؇���X�?             5@       ������������������������       �                     0@        �       �                 ��T?@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                  �>@xȂq2�?m             e@       �       �                    �?�0up[��?Y             a@        �       �                    �?8����?             7@       �       �                    �?���N8�?             5@       �       �                    �?�t����?             1@        �       �                 ���<@�����H�?             "@       ������������������������       �                     @        �       �                 X��E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @      �?              @        ������������������������       �                      @        �       �                 03�-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                     �?>A�F<�?I            �\@        �       �                 03:@l��[B��?             =@        ������������������������       �                     @        �       �                   �J@
j*D>�?             :@       �       �                 `f�;@�����?	             3@       �       �                 03k:@ףp=
�?             $@        ������������������������       �                     �?        �       �                 X�lC@�����H�?             "@        �       �                 �|�<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 X��B@X�<ݚ�?             "@       �       �                   @>@�q�q�?             @       �       �                 �|Y=@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `fF<@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?p��@���?9            @U@       �       �                    �?\#r��?*            �N@       �       �                     @ܷ��?��?(             M@       �       �                   �@@�ʈD��?            �E@       �       �                    5@ ��WV�?             :@        �       �                    &@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     6@        �       �                   @A@@�0�!��?
             1@        ������������������������       ����Q��?             @        ������������������������       �                     (@        �       �                 `�X#@�r����?             .@        �       �                    =@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             (@        ������������������������       �                     @        ������������������������       �                     8@        �       �                 �D B@      �?             @@        �       �                    �?      �?             0@        ������������������������       �                     @        �       �                 �|�<@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     0@        �                          @��U/��?F            �\@       �       �                    �?Ҿ ؞��?C            �[@       �       �                    "@0�)AU��?#            �L@        ������������������������       �                     �?        ������������������������       �        "             L@        �       �                    �?X�<ݚ�?              K@        �       �                    �?� �	��?             9@       �       �                    �?      �?             2@        �       �                 �|Y<@և���X�?             @       �       �                   �9@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �H@�eP*L��?             &@       �       �                   �5@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                 ��UO@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �                          �?J�8���?             =@        �                             @�����H�?             "@        ������������������������       �                     @                              �|�>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                  �?�G�z��?             4@                                �?      �?             2@        ������������������������       �                     �?                                 �?��.k���?             1@                               �E@և���X�?
             ,@       	                         7@      �?              @        
                      �̔Y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������C�B���?�x�z���?��؉���?ى�؉��?vb'vb'�?�N��N��?�������?�������?      �?      �?              �?^Cy�5�?(������?      �?        �?�?              �?      �?        r�q��?�q�q�?9��8���?�8��8��?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?        �������?�������?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?      �?                      �?              �?�؉�؉�?;�;��?�������?�������?333333�?�������?      �?      �?      �?                      �?      �?        �������?�������?z��y���?�a�a�?]t�E]�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?�0�9�a�?��g<�?<<<<<<�?�?      �?        /�袋.�?F]t�E�?              �?�������?�������?�k(���?(�����?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        9��8���?r�qǡ?�Cc}h��?9/���?      �?        wwwwww�?�?�؉�؉�?;�;��?      �?              �?      �?      �?                      �?      �?        ӛ���7�?d!Y�B�?      �?        }�'}�'�?l�l��?      �?      �?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?        	P� 	�?�_�����?�ڑ@;�?��K�~��?�q�q�?r�q��?�?wwwwww�?t�E]t�?]t�E�?      �?      �?              �?      �?              �?        (�����?�k(���?�������?333333�?              �?      �?                      �?UUUUUU�?UUUUUU�?6�'K`�?�d	l�O�?�7��Mo�?���,d�?'u_[�?[4���?F]t�E�?]t�E�?|���?>����?      �?      �?�a�a�?��y��y�?              �?      �?      �?�$I�$I�?n۶m۶�?              �?      �?                      �?              �?      �?        F]t�E�?/�袋.�?      �?      �?              �?      �?        �q�q�?�q�q�?UUUUUU�?�������?              �?      �?                      �?              �?]t�E�?t�E]t�?�������?ZZZZZZ�?              �?ى�؉��?�؉�؉�?      �?              �?      �?      �?                      �?      �?      �?t�E]t�?F]t�E�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?ZZZZZZ�?�������?              �?�������?�?      �?                      �?      �?        (b6�5�?aw&��+�?      �?      �?�$I�$I�?۶m۶m�?              �?333333�?�������?      �?                      �?      �?        3�E��?��1G���?��!��u�?�uy)�?d!Y�B�?8��Moz�?�a�a�?��y��y�?�������?�������?�q�q�?�q�q�?      �?              �?      �?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?������?Cy�5��?GX�i���?���=��?      �?        ;�;��?b'vb'v�?^Cy�5�?Q^Cy��?�������?�������?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?r�q��?�q�q�?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?              �?      �?        �m۶m��?�$I�$I�?      �?                      �?�������?�?��:��?XG��).�?��=���?a���{�?A_���?�}A_з?O��N���?;�;��?      �?      �?      �?      �?      �?              �?        ZZZZZZ�?�������?�������?333333�?      �?        �������?�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?              �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        g1��t�?Lg1��t�?��2���?q��$�?p�}��?��Gp�?      �?                      �?r�q��?�q�q�?)\���(�?�Q����?      �?      �?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?        t�E]t�?]t�E�?�$I�$I�?�m۶m��?      �?                      �?      �?        �$I�$I�?�m۶m��?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �rO#,��?|a���?�q�q�?�q�q�?      �?              �?      �?      �?                      �?�������?�������?      �?      �?      �?        �?�������?�$I�$I�?۶m۶m�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJL�OhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       n                     @�E	�rQ�?�           8�@               K                    �?�l�7B��?�            0r@                                  �?�a1���?�            �f@                                  �H@�nkK�?0            @Q@       ������������������������       �        '             K@                                    �?z�G�z�?	             .@                                  �?      �?              @                               ,w�U@r�q��?             @       	       
                 ���;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                   L@����X�?             @       ������������������������       �                     @        ������������������������       �                      @                                 ��$:@L�}�:G�?P            �\@                                    �?�:�]��?#            �I@        ������������������������       �                     @                                   5@dP-���?             �G@                                  �1@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                  �)@ �#�Ѵ�?            �E@        ������������������������       �                     ,@                                �|�=@ 	��p�?             =@                                   �?8�Z$���?             *@        ������������������������       �                     �?                                �|�<@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     0@        !       J                     �?p�EG/��?-            �O@       "       3                    �?���@M^�?,             O@        #       2                 �̾w@X�Cc�?             <@       $       1                   �F@ �o_��?             9@       %       0                 Ъb@��S���?             .@       &       /                 `��I@��
ц��?
             *@       '       .                    C@�eP*L��?             &@       (       -                  Y>@�q�q�?             "@       )       ,                 ���<@      �?             @        *       +                   @@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        4       I                    �?j���� �?             A@       5       >                   �F@4���C�?            �@@        6       =                   `@@X�Cc�?             ,@       7       <                 �|�?@ףp=
�?             $@       8       ;                 `fF<@z�G�z�?             @        9       :                 �|�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ?       H                    R@�d�����?             3@       @       G                  i?@@�0�!��?
             1@       A       F                    K@�z�G��?             $@       B       C                 `f�;@���Q��?             @        ������������������������       �                      @        D       E                   �=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        L       M                    �?ܧ��1�??             [@       ������������������������       �        #             P@        N       m                    �?v�X��?             F@       O       \                    <@�4F����?            �D@        P       Q                    �?�	j*D�?
             *@        ������������������������       �                     @        R       W                    �?���Q��?             $@        S       V                     �?      �?             @        T       U                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        X       Y                    �?r�q��?             @        ������������������������       �                     @        Z       [                   @9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ]       ^                   �>@؇���X�?             <@        ������������������������       �                     @        _       l                     �?r�q��?             8@       `       a                    A@"pc�
�?             6@        ������������������������       �                     �?        b       c                   �B@؇���X�?
             5@        ������������������������       �                     @        d       k                    �?@�0�!��?	             1@       e       f                 Ј�U@      �?             0@        ������������������������       �                     &@        g       j                    �?���Q��?             @       h       i                 @�pX@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        o       v                    @���L��?           @z@        p       q                    �?�<ݚ�?             2@        ������������������������       �                     "@        r       s                     @X�<ݚ�?             "@        ������������������������       �                     @        t       u                 ��T?@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        w       �                    �?z��h���?            y@        x       �                   �"@4���6��?I            @[@        y       �                 �̌@&^�)b�?            �E@       z                           �?��� ��?             ?@       {       |                 ���@�X�<ݺ?             2@        ������������������������       �                     @        }       ~                    �?�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                 ��@�θ�?	             *@       �       �                 �|�9@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?              @       �       �                   �7@r�q��?             @        ������������������������       �                     @        �       �                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �4@�q�q�?	             (@        ������������������������       �                     @        �       �                 �?�@և���X�?             @        ������������������������       �                     �?        �       �                    �?      �?             @       �       �                    9@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    @r٣����?*            �P@       �       �                    �?�c�Α�?$             M@        �       �                    �?��
ц��?             :@        ������������������������       �                     @        �       �                 ��Y.@�û��|�?             7@        �       �                 ���*@�θ�?             *@       �       �                 Ь�#@�q�q�?             "@        ������������������������       �                     @        �       �                 �[$@      �?             @        ������������������������       �                      @        �       �                 ��&@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�7@���Q��?             $@        ������������������������       �                      @        �       �                 �|Y>@      �?              @        ������������������������       �                     @        �       �                 03�1@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    @      �?             @@       �       �                   �*@$�q-�?             :@        �       �                   �&@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     6@        �       �                   @C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �                         @@@�y��>�?�            Pr@       �       �                    �?@�r-��?�            �m@        �       �                    �?�z�G��?             >@       �       �                    �?8^s]e�?             =@       �       �                 �|Y=@��+7��?             7@       �       �                    5@��
ц��?             *@        ������������������������       �                     @        �       �                    �?�q�q�?             "@       �       �                   @@      �?              @       �       �                 ���@���Q��?             @       �       �                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 �|Y7@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �                       �T�I@^���'�?�            �i@       �       �                    �?T�Ü&�?~            �h@        �       �                  ��@�MI8d�?            �B@        ������������������������       �                     "@        �       �                    �?d}h���?             <@       �       �                 �|Y=@�z�G��?
             4@        ������������������������       �                      @        �       �                 ��(@�<ݚ�?	             2@       ������������������������       �      �?             0@        ������������������������       �                      @        ������������������������       �                      @        �       �                    $@�����H�?i            @d@        �       �                    @���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �>@P��-�?d            �c@       �       �                 �?�@�L���?]            �b@        �       �                   �7@��?^�k�?-            �Q@        ������������������������       �                     6@        �       �                 ���@ �q�q�?             H@        �       �                    �?      �?             @       �       �                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?`���i��?             F@       �       �                 �|Y=@ qP��B�?            �E@        ������������������������       �                     6@        �       �                  sW@���N8�?             5@        �       �                 pf�@؇���X�?             @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �        	             ,@        ������������������������       �                     �?        �       �                   �4@�ݜ�?0            �S@        �       �                 ��Y @r֛w���?             ?@        �       �                   �2@�q�q�?             (@        ������������������������       �                      @        �       �                 @3�@���Q��?             $@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �3@և���X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     3@        �       �                 ��) @`�q�0ܴ?            �G@        ������������������������       �                     8@        �       �                   �:@���}<S�?             7@        ������������������������       �                      @        �       �                   �;@�r����?
             .@        ������������������������       �                     �?        �       �                 pf� @@4և���?	             ,@        ������������������������       �                     �?        ������������������������       �                     *@        �                       ��I @�q�q�?             "@                                �?@և���X�?             @        ������������������������       �                      @                              �?�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @                              p�O@և���X�?             @             
                �|�>@      �?             @             	                   ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                              �?�@0�)AU��?$            �L@        ������������������������       �                     ?@                                 �? ��WV�?             :@                                �?P���Q�?             4@                             @3�@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     �?        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������JP���?7j_Q��?�X){�+�?�Sk���?�/���?�7�v���?d!Y�B�?�Mozӛ�?              �?�������?�������?      �?      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�$I�$I�?�m۶m��?              �?      �?        �}���?~��G�?}}}}}}�?�?      �?        �����F�?W�+�ɵ?      �?      �?      �?                      �?�/����?�}A_Ч?      �?        ������?�{a���?;�;��?;�;��?      �?        �������?UUUUUU�?      �?                      �?      �?        �4M�4M�?Y�eY�e�?�s�9��?�c�1��?%I�$I��?�m۶m��?
ףp=
�?�Q����?�?�������?�؉�؉�?�;�;�?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?                      �?              �?      �?                      �?              �?      �?              �?                      �?�������?ZZZZZZ�?m��&�l�?'�l��&�?�m۶m��?%I�$I��?�������?�������?�������?�������?      �?      �?              �?      �?                      �?              �?      �?        Cy�5��?y�5���?ZZZZZZ�?�������?ffffff�?333333�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?      �?                      �?�%���^�?	�%����?              �?�.�袋�?颋.���?ە�]���?KԮD�J�?;�;��?vb'vb'�?              �?�������?333333�?      �?      �?      �?      �?      �?                      �?      �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?/�袋.�?F]t�E�?              �?۶m۶m�?�$I�$I�?      �?        ZZZZZZ�?�������?      �?      �?      �?        333333�?�������?      �?      �?              �?      �?                      �?              �?      �?              �?        ��:��:�?_�_��?�q�q�?9��8���?              �?�q�q�?r�q��?              �?�������?�������?      �?                      �?��C���?t��2�?q=��?߅����?�}A_��?���/��?�B!��?�{����?�q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?              �?      �?        �؉�؉�?ى�؉��?�������?333333�?              �?      �?              �?      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?�$I�$I�?۶m۶m�?      �?              �?      �?�������?333333�?      �?                      �?      �?        >���>�?|���?5�rO#,�?�{a���?�;�;�?�؉�؉�?              �?8��Moz�?��,d!�?ى�؉��?�؉�؉�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        �������?333333�?      �?              �?      �?              �?�������?333333�?              �?      �?              �?      �?�؉�؉�?;�;��?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ������?���E�)�?'u_�?��c+���?ffffff�?333333�?|a���?	�=����?zӛ����?Y�B��?�;�;�?�؉�؉�?      �?        UUUUUU�?UUUUUU�?      �?      �?�������?333333�?      �?      �?              �?      �?              �?                      �?      �?              �?              �?      �?      �?                      �?      �?        Y�'�J��?��`����?�xN%$�?�8���߾?��L���?L�Ϻ��?      �?        I�$I�$�?۶m۶m�?ffffff�?333333�?              �?9��8���?�q�q�?      �?      �?      �?              �?        �q�q�?�q�q�?�������?333333�?              �?      �?        6��(S��?R��fu�?}���g�?L�Ϻ��?_�_��?�A�A�?      �?        �������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        F]t�E�?F]t�E�?��}A�?�}A_З?      �?        ��y��y�?�a�a�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?        \��[���?�i�i�?���{��?�B!��?UUUUUU�?UUUUUU�?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?        ��F}g��?W�+�ɥ?      �?        ӛ���7�?d!Y�B�?      �?        �������?�?              �?n۶m۶�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?�������?�������?      �?              �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?                      �?      �?        ��Gp�?p�}��?      �?        O��N���?;�;��?ffffff�?�������?�5��P�?(�����?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��lhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       J                     �?>AU`�z�?�           8�@               	                    �?�û��|�?v             g@                                   !@�g<a�?/            @S@        ������������������������       �                     �?                                83A@�"w����?.             S@                                ���;@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        *            �Q@        
       I                   �J@�E1���?G            �Z@                                 �;@h�|�`�?9            �U@                                   9@������?	             .@                                  �?      �?              @                               ���Q@�q�q�?             @        ������������������������       �                      @                                  �4@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               H                 p�w@"` Y��?0            �Q@              1                  �>@.Lj���?.             Q@               0                    �?l��[B��?             =@                                  �?
j*D>�?             :@                                �|�=@      �?             @                               �ܵ<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                03:@8�A�0��?             6@        ������������������������       �                     @                !                 03k:@     ��?
             0@        ������������������������       �                     @        "       /                   @>@�θ�?	             *@       #       ,                 `fF<@�z�G��?             $@       $       '                 �|�?@����X�?             @        %       &                 �|�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        (       )                   �C@z�G�z�?             @        ������������������������       �                     @        *       +                    H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        -       .                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        2       9                    �?x�����?            �C@       3       8                    �?���N8�?             5@        4       7                 `f�A@؇���X�?             @        5       6                  �>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        :       ;                   �B@b�2�tk�?             2@        ������������������������       �                     @        <       C                    �?��
ц��?	             *@       =       B                   �H@�q�q�?             @       >       A                    �?      �?             @       ?       @                 �U�T@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        D       E                   �E@����X�?             @        ������������������������       �                     @        F       G                   �G@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@        K       �                    �?�[Yqf��?O           x�@       L       S                    /@�3�E���?            z@        M       N                    �?r�q��?             (@        ������������������������       �                     @        O       P                 �&�)@����X�?             @        ������������������������       �                     @        Q       R                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        T       �                    �?�zӝ���?           @y@        U       \                 ��@�ț��*�??            �W@        V       [                 P�@�}�+r��?             3@        W       X                    �?z�G�z�?             @        ������������������������       �                      @        Y       Z                 �|Y:@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             ,@        ]       r                    �?|�i���?1             S@       ^       _                    �?8����?             G@        ������������������������       �                     @        `       e                   �9@#z�i��?            �D@        a       b                 @�"@      �?             (@       ������������������������       �                     @        c       d                    4@      �?             @        ������������������������       �                     @        ������������������������       �                     @        f       k                     @д>��C�?             =@       g       h                   �B@�}�+r��?             3@       ������������������������       �                     &@        i       j                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        l       m                    ;@���Q��?             $@        ������������������������       �                     @        n       o                 ��� @z�G�z�?             @        ������������������������       �                     @        p       q                  SE"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        s       t                 P�@�z�G��?             >@        ������������������������       �                     @        u       v                 ��'@�q�q�?             ;@        ������������������������       �                      @        w       ~                     @ �o_��?             9@       x       y                 ��m1@�	j*D�?	             *@        ������������������������       �                      @        z       {                   �7@���|���?             &@        ������������������������       �                      @        |       }                   �E@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @               �                 �|�;@      �?             (@        ������������������������       �                      @        �       �                    �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    A@,���j�?�            Ps@       �       �                    �?�E�X̚�?�            �o@       �       �                     @��[��?�            �k@        �       �                    �?R���Q�?             D@        ������������������������       �                     @        �       �                   �@@�MI8d�?            �B@       �       �                 �|�=@�t����?             A@       �       �                   �3@PN��T'�?             ;@       �       �                   �(@"pc�
�?             6@        �       �                    &@؇���X�?             ,@       �       �                    5@"pc�
�?             &@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|Y;@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                   �7@�1j�P�?t            �f@        �       �                    �?h㱪��?"            �K@        ������������������������       �                      @        �       �                 @3�@�&=�w��?!            �J@       ������������������������       �                     <@        �       �                 0S5 @HP�s��?             9@        �       �                   �3@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     5@        �       �                 ��) @�ŇG+��?R            �_@       �       �                    �?�>����?G             [@        �       �                 ���@��-�=��?            �C@        ������������������������       �                     $@        �       �                 ���@\-��p�?             =@        �       �                 �|�=@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                 P�J@�8��8��?             8@       �       �                  ��@�r����?             .@        ������������������������       �                     @        �       �                 �|Y=@z�G�z�?             $@        ������������������������       �                     �?        ������������������������       ������H�?             "@        ������������������������       �                     "@        �       �                 �?$@p��%���?-            @Q@        �       �                 �&b@؇���X�?             5@        ������������������������       �                     "@        �       �                 ���@      �?	             (@        ������������������������       �                      @        �       �                 �|Y;@ףp=
�?             $@        ������������������������       �                     @        �       �                 �|Y>@r�q��?             @       �       �                 pf�@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �?�@@��8��?!             H@       ������������������������       �                     :@        �       �                    ?@���7�?             6@       ������������������������       �                     1@        �       �                 @3�@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                 �!�A@      �?             2@       �       �                    ?@���Q��?	             .@       �       �                    (@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    6@      �?             @@       ������������������������       �                     8@        �       �                     @      �?              @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�@�h����?"             L@        �       �                    �?h�����?             <@        ������������������������       �                     $@        �       �                   �D@�X�<ݺ?
             2@        �       �                   @C@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     <@        �                          �;@�f��`��?G            �[@       �       �                    !@�	j*D�?+            @P@       �       �                     @"pc�
�?            �@@        ������������������������       �                     &@        �       �                 03�9@���!pc�?             6@       �       �                    �?�8��8��?	             (@        ������������������������       �                     @        �       �                    @�����H�?             "@        �       �                 pf�0@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             $@        ������������������������       �                     �?        �       �                    @X�<ݚ�?             "@        ������������������������       �                     @        �       �                 ��T?@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?     ��?             @@       �       �                    �?8����?             7@       �       �                    �?�����H�?             2@       �       �                     @"pc�
�?             &@        ������������������������       �                     @        �       �                    +@�q�q�?             @        ������������������������       �                     �?        �       �                   �6@z�G�z�?             @       �       �                 ��'@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `f2@�<ݚ�?             "@        �       �                 `ff+@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                 �?���j��?             G@                                �?����"�?             =@                              �|Y>@      �?              @       ������������������������       �                     @        ������������������������       �                      @                                 �?���N8�?             5@        ������������������������       �                     �?              	                032@z�G�z�?             4@        ������������������������       �                      @        
                         �?�q�q�?	             (@                             `fV6@      �?              @        ������������������������       �                      @                                �>@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                 @�t����?
             1@        ������������������������       �                      @                                 �?�<ݚ�?             "@        ������������������������       �                     @                                 �?���Q��?             @                                 @�q�q�?             @        ������������������������       �                     �?                              pf�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?��,d!�?8��Moz�?�cj`?���8+�?      �?        (�����?Cy�5��?UUUUUU�?�������?              �?      �?                      �?Q�@��?]���~!�?��#�;�?⎸#��?�?wwwwww�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?�V�H�?��RO�o�?------�?�������?GX�i���?���=��?;�;��?b'vb'v�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        /�袋.�?颋.���?      �?              �?      �?              �?�؉�؉�?ى�؉��?333333�?ffffff�?�$I�$I�?�m۶m��?      �?      �?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ��o��o�?�A�A�?��y��y�?�a�a�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �8��8��?9��8���?      �?        �؉�؉�?�;�;�?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?              �?      �?        �5_���?)�A��(�?;�;��?ى�؉��?UUUUUU�?�������?              �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?�(0��<�?�]?[��?�a�+�?�~�-q��?(�����?�5��P�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�5��P^�?�5��P�?8��Moz�?d!Y�B�?              �?ە�]���?�+Q��?      �?      �?      �?              �?      �?              �?      �?        |a���?a���{�?(�����?�5��P�?              �?      �?      �?      �?                      �?�������?333333�?              �?�������?�������?      �?              �?      �?              �?      �?        333333�?ffffff�?              �?UUUUUU�?UUUUUU�?      �?        �Q����?
ףp=
�?;�;��?vb'vb'�?              �?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?              �?      �?              �?      �?      �?        �������?�������?      �?                      �?<�o�14�?#>�Tr^�?�5g"��?��R��N�?�Ma�Ma�?�����?333333�?333333�?      �?        ��L���?L�Ϻ��?<<<<<<�?�?&���^B�?h/�����?/�袋.�?F]t�E�?۶m۶m�?�$I�$I�?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?              �?              �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?������?�8xߺ?־a���?��)A��?      �?        tHM0���?�x+�R�?      �?        q=
ףp�?{�G�z�?      �?      �?              �?      �?              �?        캮뺮�?QEQE�?�Kh/��?h/�����?}˷|˷�?�A�A�?      �?        a����?�{a���?333333�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?�������?�?      �?        �������?�������?              �?�q�q�?�q�q�?      �?        �g��%�?ہ�v`��?۶m۶m�?�$I�$I�?      �?              �?      �?              �?�������?�������?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?        �.�袋�?F]t�E�?      �?        �������?�������?      �?      �?      �?              �?      �?333333�?�������?]t�E�?t�E]t�?              �?      �?              �?                      �?      �?      �?      �?              �?      �?      �?              �?      �?      �?                      �?۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?      �?        ��8��8�?�q�q�?      �?      �?      �?                      �?      �?              �?        �蕱���?�5'���?;�;��?vb'vb'�?F]t�E�?/�袋.�?              �?t�E]t�?F]t�E�?UUUUUU�?UUUUUU�?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?        �q�q�?r�q��?      �?        UUUUUU�?�������?      �?                      �?      �?      �?8��Moz�?d!Y�B�?�q�q�?�q�q�?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        9��8���?�q�q�?333333�?�������?      �?                      �?      �?        ozӛ���?!Y�B�?	�=����?�i��F�?      �?      �?              �?      �?        �a�a�?��y��y�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        <<<<<<�?�?      �?        9��8���?�q�q�?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�-#hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM=hjh))��}�(h,h/h0M=��h2h3h4hph<�h=Kub������       �                     @ʡ�;S��?�           8�@               a                  x#J@�F�i*��?�            �s@                                  @�
[���?�            `i@        ������������������������       �                      @               "                    �??����?            `h@               !                    �?L������?+            @R@              
                 `f�)@�Z��L��?)            �Q@               	                   �J@���7�?	             6@       ������������������������       �                     5@        ������������������������       �                     �?                                    �?؇���X�?             �H@                                   �?؇���X�?             @                                  �?r�q��?             @                                hލC@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                   �?؇���X�?             E@                                  �<@�LQ�1	�?             7@                                  �+@�q�q�?             "@                                   5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@                                   �E@�S����?             3@                                  6@�����H�?             2@                                ��m1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �                     �?        ������������������������       �                      @        #       P                    �?`��:�?T            �^@       $       -                    �?�v�G���?F            �Y@        %       ,                    �?      �?              @       &       +                   �A@և���X�?             @       '       (                  `6@���Q��?             @        ������������������������       �                     �?        )       *                 X��E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        .       =                     �?fGk�T�??            �W@        /       <                    �?f���M�?             ?@       0       1                 �|�<@����"�?             =@        ������������������������       �                      @        2       ;                  i?@�q�q�?             ;@       3       4                    D@��.k���?             1@        ������������������������       �                     @        5       6                   �G@�n_Y�K�?             *@        ������������������������       �                     @        7       :                 `fF<@����X�?             @       8       9                   �K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             $@        ������������������������       �                      @        >       O                    �?     �?(             P@       ?       N                   �*@�IєX�?#            �I@       @       E                 `f�)@�L���?            �B@        A       D                    &@��S�ۿ?             .@       B       C                    5@$�q-�?	             *@        ������������������������       �      �?             @        ������������������������       �                     "@        ������������������������       �                      @        F       G                 �|�<@�C��2(�?             6@        ������������������������       �                     "@        H       I                 �|�=@8�Z$���?
             *@        ������������������������       �                     �?        J       M                   �A@�8��8��?	             (@        K       L                    @@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     *@        Q       V                    :@p�ݯ��?             3@        R       U                    �?և���X�?             @       S       T                    *@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        W       ^                    �?      �?             (@       X       Y                    �?�����H�?             "@        ������������������������       �                      @        Z       [                   P@@؇���X�?             @        ������������������������       �                     @        \       ]                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        _       `                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        b       �                  "�b@�*�Lk�?F            @\@       c       n                    �?д>��C�?7            �U@        d       e                    �?�˹�m��?             C@       ������������������������       �                     >@        f       m                 ��!T@      �?              @       g       l                     �?      �?             @       h       i                   �9@�q�q�?             @        ������������������������       �                     �?        j       k                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        o       �                   �P@ \� ���?             �H@       p       �                 �\@��[�p�?            �G@       q       �                   �I@      �?             D@       r       y                    �?     ��?             @@        s       t                 p"�X@�d�����?             3@       ������������������������       �                     &@        u       v                    �?      �?              @        ������������������������       �                     @        w       x                    F@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        z       �                 03sP@�n_Y�K�?             *@       {       �                 03�O@���!pc�?
             &@       |       }                   �A@      �?              @        ������������������������       �                     @        ~                        `�iJ@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?��
ц��?             :@       �       �                    !@      �?	             0@        ������������������������       �                     @        ������������������������       �                     $@        �       �                 03c@z�G�z�?             $@        ������������������������       �                     �?        �       �                    �?�����H�?             "@       �       �                 �̾w@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���@�6�W�?�            �x@        ������������������������       �                     <@        �       �                    �?�$Jd��?�            �v@        �       �                 `v�6@�AMĹ�?C             [@       �       �                    �?(Q��h�?3            @T@        �       �                    �?��Sݭg�?            �C@        �       �                    �?b�2�tk�?
             2@        ������������������������       �                     @        �       �                    �?��
ц��?             *@       �       �                 `�@1@      �?             (@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|Y8@؇���X�?             5@        ������������������������       �                     @        �       �                    �?@�0�!��?             1@       �       �                    �?��S�ۿ?             .@       �       �                  ��@$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                      @        �       �                 ��Y1@�D����?             E@       �       �                 `f�%@��%��?            �B@       �       �                    @d��0u��?             >@       �       �                    �?J�8���?             =@       �       �                   �5@�q�q�?             ;@        �       �                    �?�<ݚ�?             "@       �       �                 @�"@�q�q�?             @       �       �                   �4@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�����H�?
             2@       �       �                 ���@      �?	             0@        �       �                 �|Y:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 pf� @@4և���?             ,@       �       �                    ;@؇���X�?             @        �       �                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �;@؇���X�?             @        ������������������������       �                     @        �       �                 �|�<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�����H�?             ;@        ������������������������       �                      @        �       �                 ��T?@`2U0*��?             9@       ������������������������       �                     5@        �       �                    @      �?             @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �                       ��M%@+����?�            0p@       �                          �?�A����?m             g@       �       �                 ��@t���s��?i             f@        ������������������������       �                     �?        �       �                    �?L���#��?h             f@        �       �                 ���@8�Z$���?             :@        ������������������������       �                     @        �       �                 �� @���y4F�?
             3@       �       �                   �5@����X�?	             ,@        ������������������������       �                     �?        �       �                   �<@�θ�?             *@        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             "@        ������������������������       �                     �?        �       �                   @@      �?              @       ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    :@ףp=
�?X            �b@        �       �                    �?P���Q�?!             N@        ������������������������       �                      @        �       �                 @3�@�8���?              M@        ������������������������       �                     9@        �       �                 pf� @�C��2(�?            �@@        �       �                   �3@@�0�!��?             1@        �       �                   �1@և���X�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �        	             0@        �                       @Q!@�r����?7            �V@       �       �                   �>@�����?.            �R@       �       �                    �? �#�Ѵ�?            �E@        �       �                 �Y�@r�q��?             @        ������������������������       �                     �?        �       �                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?$@�?�|�?            �B@        �       �                 ��@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     >@        �       �                   �?@�חF�P�?             ?@        ������������������������       �                     @                                  �?@4և���?             <@        ������������������������       �                     @                                �B@HP�s��?             9@        ������������������������       �                     &@                                �D@؇���X�?             ,@        ������������������������       ����Q��?             @        ������������������������       �                     "@              
                0S%"@     ��?	             0@              	                �|Y<@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                              ���"@"pc�
�?             &@        ������������������������       �                     �?                                �<@z�G�z�?             $@        ������������������������       �                     @                              �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                 �?����X�?             @                                �?���Q��?             @        ������������������������       �                      @                              P�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                              0S�*@�+e�X�?-            �R@        ������������������������       �                     @              <                  @@@�㙢�c�?*            @Q@             !                   �?���y4F�?$            �L@                                  �?r�q��?             @                             �0@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        "      9                �|�>@L紂P�?!            �I@       #      2                   �?8��8���?             H@       $      +                   �?��(\���?             D@       %      *                   �?�>����?             ;@        &      '                  `3@      �?             @        ������������������������       �                     �?        (      )                03�7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        ,      -                   !@$�q-�?
             *@       ������������������������       �                     $@        .      1                   @�q�q�?             @       /      0                   +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        3      8                    @      �?              @        4      5                �̌4@�q�q�?             @        ������������������������       �                     �?        6      7                   +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        :      ;                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        �*       h�h))��}�(h,h/h0M=KK��h2h3h4hVh<�h=Kub������������N���I5�?d�~`l��?��JG��?
�Z܄�?б�n��?�_�"�?      �?        QeQe�?]�5]�5�?����?�Ǐ?~�?��Vؼ?���.�d�?F]t�E�?�.�袋�?              �?      �?        �$I�$I�?۶m۶m�?�$I�$I�?۶m۶m�?UUUUUU�?�������?      �?      �?      �?                      �?              �?              �?�$I�$I�?۶m۶m�?Y�B��?��Moz��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?^Cy�5�?(������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?*.�u��?XG��).�?C���?��O �?      �?      �?�$I�$I�?۶m۶m�?�������?333333�?      �?              �?      �?              �?      �?              �?              �?        ��c�H�?�-q����?��RJ)��?��Zk���?	�=����?�i��F�?              �?UUUUUU�?UUUUUU�?�?�������?              �?;�;��?ى�؉��?      �?        �$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?              �?             ��?      �?�?�?}���g�?L�Ϻ��?�������?�?�؉�؉�?;�;��?      �?      �?      �?              �?        ]t�E�?F]t�E�?      �?        ;�;��?;�;��?              �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?              �?              �?        ^Cy�5�?Cy�5��?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?              �?      �?�q�q�?�q�q�?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ��M�l�?�|٠��?|a���?a���{�?^Cy�5�?��P^Cy�?              �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?և���X�?
^N��)�?m�w6�;�?�
br1�?      �?      �?      �?      �?y�5���?Cy�5��?              �?      �?      �?      �?              �?      �?              �?      �?        ى�؉��?;�;��?t�E]t�?F]t�E�?      �?      �?              �?333333�?�������?              �?      �?                      �?      �?                      �?              �?      �?        �;�;�?�؉�؉�?      �?      �?      �?                      �?�������?�������?              �?�q�q�?�q�q�?�������?�������?      �?                      �?      �?        ��$5��?�;l+��?      �?        c�Zb=�?�sF�v
�?���^B{�?��^B{	�?������?x�5?,�?�i�i�?�|˷|��?9��8���?�8��8��?              �?�;�;�?�؉�؉�?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?�������?ZZZZZZ�?�?�������?;�;��?�؉�؉�?      �?                      �?              �?      �?        �0�0�?z��y���?���L�?}���g�?DDDDDD�?wwwwww�?�rO#,��?|a���?UUUUUU�?UUUUUU�?�q�q�?9��8���?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�q�q�?�q�q�?      �?      �?      �?      �?              �?      �?        n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?              �?              �?      �?              �?      �?                      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?�q�q�?              �?���Q��?{�G�z�?      �?              �?      �?      �?      �?      �?                      �?      �?        �o���?K<A���?C���,�?�Mozӛ�?3��Yb�?k��2�?              �?�.�袋�?��.�袻?;�;��?;�;��?      �?        6��P^C�?(������?�m۶m��?�$I�$I�?              �?ى�؉��?�؉�؉�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?333333�?�������?      �?              �?        �������?�������?ffffff�?�������?      �?        j��FX�?a���{�?      �?        ]t�E�?F]t�E�?ZZZZZZ�?�������?�$I�$I�?۶m۶m�?�������?�������?              �?      �?              �?        �������?�?�Ϻ���?v�)�Y7�?�/����?�}A_Ч?�������?UUUUUU�?      �?        �������?�������?              �?      �?        *�Y7�"�?к����?۶m۶m�?�$I�$I�?      �?              �?      �?      �?        �Zk����?��RJ)��?              �?n۶m۶�?�$I�$I�?      �?        q=
ףp�?{�G�z�?      �?        ۶m۶m�?�$I�$I�?333333�?�������?      �?              �?      �?�������?333333�?              �?      �?        /�袋.�?F]t�E�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        R���Q�?���Q��?              �?�7��Mo�?d!Y�B�?6��P^C�?(������?UUUUUU�?�������?      �?      �?      �?                      �?              �?�������?�������?�������?�������?�������?333333�?�Kh/��?h/�����?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ5�;5hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMChjh))��}�(h,h/h0MC��h2h3h4hph<�h=Kub������       �                    �?�3)0�F�?�           8�@              �                    �?^����?T           h�@              �                 03S@��iŪ��?           �x@                               ���@�KaW\�?�            �w@        ������������������������       �                     9@               w                   `@@h &A�l�?�            Pv@              l                   �?@�ĚpF�?�            �o@                                  �?<�yr��?�            �n@        	       
                    �?L紂P�?             �I@        ������������������������       �                     9@                                �|�=@R�}e�.�?             :@                               �|Y=@�X����?             6@                                 �7@      �?             4@                                   @     ��?             0@        ������������������������       �                     @                                pf�@�θ�?             *@        ������������������������       �                     @                                   '@      �?              @        ������������������������       �                     �?                                 �#@և���X�?             @                                  4@���Q��?             @        ������������������������       �                      @                                �̜!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                  �<@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                '                 �Y�@ʨ����?~             h@        !       &                   �8@�\��N��?
             3@        "       #                   �6@�C��2(�?             &@        ������������������������       �                      @        $       %                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        (       a                 `fF:@\-��p�?t            �e@       )       *                 ���@,I�e���?e            �b@        ������������������������       �                     3@        +       @                   �<@��U�=��?Y            �`@        ,       -                 @3�@`Jj��?,             O@        ������������������������       �                     7@        .       ;                   �3@��-�=��?            �C@        /       0                 pf� @�S����?             3@        ������������������������       �                      @        1       2                    �?�IєX�?
             1@        ������������������������       �                      @        3       4                   �2@��S�ۿ?	             .@       ������������������������       �                     $@        5       6                 ���$@z�G�z�?             @        ������������������������       �                      @        7       :                     @�q�q�?             @       8       9                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        <       =                 ��q1@P���Q�?             4@       ������������������������       �                     2@        >       ?                 ��d6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        A       D                    �?z��R[�?-            �Q@        B       C                 �|Y=@      �?              @        ������������������������       �                     @        ������������������������       �                     @        E       N                 ��) @�חF�P�?)             O@       F       G                    �?�L���?            �B@        ������������������������       �z�G�z�?             $@        H       M                 �|�=@ 7���B�?             ;@       I       J                 �|Y=@�nkK�?             7@        ������������������������       �                     �?        K       L                  sW@���7�?             6@        ������������������������       �      �?              @        ������������������������       �                     4@        ������������������������       �                     @        O       `                   �>@ �o_��?             9@       P       Q                 `��!@�q�q�?             8@        ������������������������       �                      @        R       _                   �+@�GN�z�?             6@       S       X                     @�q�q�?	             .@       T       W                 �|�=@�q�q�?             @        U       V                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        Y       ^                 �|�=@�q�q�?             "@       Z       ]                 �|Y=@؇���X�?             @       [       \                 ���"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        b       e                   �<@8����?             7@        c       d                   �7@      �?              @        ������������������������       �                      @        ������������������������       �                     @        f       g                 �|Y=@��S�ۿ?
             .@        ������������������������       �                      @        h       k                    �?$�q-�?	             *@        i       j                 ��2>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        m       r                     @�eP*L��?             &@        n       q                    @@      �?             @       o       p                   �'@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        s       v                 d�@@և���X�?             @       t       u                 �?�@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        x       �                     @��x_F-�?B            �Y@       y       �                    �?��M���?-             Q@        z                        ���;@"pc�
�?             &@       {       |                   �J@ףp=
�?             $@       ������������������������       �                     @        }       ~                   �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��$:@�k�'7��?&            �L@        �       �                    �?(;L]n�?             >@        ������������������������       �                     @        �       �                   @A@ �q�q�?             8@        ������������������������       �      �?              @        ������������������������       �                     6@        �       �                   �J@�q�q�?             ;@       �       �                   �G@      �?             0@       �       �                   �F@�n_Y�K�?
             *@       �       �                    �?      �?              @        �       �                    C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    D@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                  Y>@�C��2(�?             &@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?г�wY;�?             A@        ������������������������       �                     @        �       �                   �C@ 7���B�?             ;@       �       �                   @C@ףp=
�?	             $@       ������������������������       �                     @        �       �                 ��	0@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �        
             ,@        �       �                     �?v ��?R             `@        �       �                    �?��Hg���?            �F@       �       �                    �?���N8�?             E@       ������������������������       �                     5@        �       �                 p"�X@�G��l��?             5@       �       �                    �?b�2�tk�?
             2@        ������������������������       �                     @        �       �                    D@���|���?             &@       �       �                 03�Q@և���X�?             @       �       �                    7@���Q��?             @        ������������������������       �                      @        �       �                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��i#[�?4             U@        �       �                 038@�q�q�?             8@       �       �                    �?      �?             0@       �       �                    3@������?             .@        ������������������������       �                     �?        �       �                     @d}h���?
             ,@        �       �                 ���2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?r�q��?             (@        �       �                  S�-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                      @        �       �                     @������?$             N@        �       �                    �? �o_��?             9@       �       �                    6@�q�q�?             8@        ������������������������       �                      @        �       �                   �7@�GN�z�?             6@        ������������������������       �                     $@        �       �                   �C@�q�q�?	             (@       �       �                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��R[s�?            �A@        �       �                 �|�;@      �?             0@       �       �                 P�@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��Y.@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    5@�}�+r��?             3@        �       �                  s�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             1@        �                       03�3@nCJ6��?u            @g@        �       �                     @8����?             G@        �       �                    �?r�q��?             (@       ������������������������       �                      @        �       �                    *@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?ҳ�wY;�?             A@       �       �                    �?�\��N��?             3@       �       �                 `�@1@���|���?             &@       �       �                    &@�z�G��?             $@        ������������������������       �                      @        �       �                 03�-@      �?              @       ������������������������       �                     @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?              @       �       �                   �2@؇���X�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 xF4!@z�G�z�?
             .@        ������������������������       �                     �?        �                          �?؇���X�?	             ,@       �                          �;@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?                                 �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @              (                ��H@�G�z��?V            �a@                                 @P�%f��?9            �V@                                 �?r٣����?            �@@       ������������������������       �                     2@        	      
                  �0@��S���?             .@        ������������������������       �                     @        ������������������������       �                      @                                 �?�KM�]�?&            �L@        ������������������������       �                     @                                 @ȵHPS!�?"             J@                                 �?      �?
             0@        ������������������������       �                     @                                 @X�<ݚ�?             "@        ������������������������       �                     @                                 �?r�q��?             @                              ��T?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @              '                   �?�X�<ݺ?             B@              &                   �?8�Z$���?             *@                                �?�<ݚ�?             "@        ������������������������       �                     @              %                   @�q�q�?             @                                  @���Q��?             @                                �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        !      "                ��T?@�q�q�?             @        ������������������������       �                     �?        #      $                ��p@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        )      B                   @��H�}�?             I@       *      A                   @8����?             G@       +      @                    �?���X�K�?            �F@       ,      3                  �B@��i#[�?             E@       -      .                   �?��2(&�?             6@        ������������������������       �                     $@        /      2                   �?      �?             (@        0      1                ��f`@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        4      5                  @C@      �?             4@        ������������������������       �                     @        6      ?                hDba@j���� �?
             1@       7      >                   �?��
ц��?             *@       8      ;                  �J@�z�G��?             $@       9      :                   F@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        <      =                  �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MCKK��h2h3h4hVh<�h=Kub������������Rl���?�[�'��?쌛�&�?�'�����?���v�?gH���?qT��I�?W��l�?      �?        �������?���?uuuuuu�?�?�h�>��?�).�u�?�������?�������?              �?�;�;�?'vb'vb�?]t�E]�?�E]t��?      �?      �?      �?      �?              �?�؉�؉�?ى�؉��?              �?      �?      �?              �?۶m۶m�?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?      �?                      �?�+���\�?�P�ݙ��?�5��P�?y�5���?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        a����?�{a���?�q˸e�?�Hs�9Ҽ?      �?        �>���?|��|�?���{��?�B!��?      �?        }˷|˷�?�A�A�?(������?^Cy�5�?              �?�?�?      �?        �������?�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        ffffff�?�������?      �?              �?      �?              �?      �?        ���?X|�W|��?      �?      �?              �?      �?        �Zk����?��RJ)��?}���g�?L�Ϻ��?�������?�������?	�%����?h/�����?�Mozӛ�?d!Y�B�?      �?        �.�袋�?F]t�E�?      �?      �?      �?              �?        
ףp=
�?�Q����?�������?�������?              �?�袋.��?]t�E�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?              �?        d!Y�B�?8��Moz�?      �?      �?      �?                      �?�������?�?      �?        �؉�؉�?;�;��?      �?      �?              �?      �?              �?        ]t�E�?t�E]t�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?۶m۶m�?�$I�$I�?333333�?�������?      �?              �?      �?              �?�������?�?�?�������?F]t�E�?/�袋.�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        -����b�?Lg1��t�?�������?�?      �?        �������?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?;�;��?ى�؉��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �?�?      �?        	�%����?h/�����?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?                      �?G�w��?qG�w��?��I��I�?؂-؂-�?��y��y�?�a�a�?              �?��y��y�?1�0��?9��8���?�8��8��?              �?]t�E]�?F]t�E�?۶m۶m�?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�a�a�?�<��<��?�������?�������?      �?      �?wwwwww�?�?              �?I�$I�$�?۶m۶m�?      �?      �?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?              �?      �?        wwwwww�?�?
ףp=
�?�Q����?�������?�������?              �?�袋.��?]t�E�?      �?        �������?�������?�$I�$I�?�m۶m��?              �?      �?              �?              �?        X|�W|��?PuPu�?      �?      �?      �?      �?              �?      �?              �?      �?      �?                      �?�5��P�?(�����?      �?      �?      �?                      �?      �?        P?���O�?X`�X�?8��Moz�?d!Y�B�?UUUUUU�?�������?              �?      �?      �?      �?                      �?�������?�������?�5��P�?y�5���?]t�E]�?F]t�E�?ffffff�?333333�?              �?      �?      �?      �?              �?      �?              �?      �?                      �?      �?      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?        �������?�������?      �?        �$I�$I�?۶m۶m�?�������?�������?              �?      �?              �?      �?      �?                      �?�������?�������?�O��O��?�`�`�?|���?>���>�?              �?�?�������?              �?      �?        �k(���?(�����?      �?        ��N��N�?�؉�؉�?      �?      �?      �?        r�q��?�q�q�?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        ��8��8�?�q�q�?;�;��?;�;��?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?              �?        
ףp=
�?{�G�z�?8��Moz�?d!Y�B�?�'}�'}�?l�l��?�<��<��?�a�a�?t�E]t�?��.���?              �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?      �?        ZZZZZZ�?�������?�;�;�?�؉�؉�?ffffff�?333333�?۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJi4�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM#hjh))��}�(h,h/h0M#��h2h3h4hph<�h=Kub������       |                     @H���I�?�           8�@               )                    �?(*Gh���?�            0s@                                  �6@4�B��?4            �R@        ������������������������       �        	             *@               $                     �?�u���?+            �N@              #                    �?�t����?%            �I@                                 @H@ �o_��?$             I@                                  C@@�0�!��?             A@       	                          �A@�+e�X�?             9@       
                           �?��2(&�?             6@                                  �?r�q��?             2@       ������������������������       �                     &@                                  �7@և���X�?             @        ������������������������       �                      @                                ��9K@���Q��?             @        ������������������������       �                     �?                                   �?      �?             @                               p�w@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@                                    �?      �?
             0@                               м�J@      �?             (@        ������������������������       �                     @                                   �?�q�q�?             "@       ������������������������       �                     @                                �UkT@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        !       "                   @J@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        %       &                    �?ףp=
�?             $@        ������������������������       �                      @        '       (                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        *       A                    �?.�����?�             m@        +       >                    :@�KM�]�?;            �W@        ,       7                   �B@&^�)b�?            �E@       -       6                   �;@ܷ��?��?             =@       .       /                   �'@�S����?             3@        ������������������������       �                     @        0       1                   �+@�θ�?	             *@        ������������������������       �                      @        2       5                    �?�C��2(�?             &@        3       4                   �9@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             $@        8       =                   @F@X�Cc�?             ,@        9       <                   �E@      �?              @       :       ;                   �C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ?       @                    @ ��WV�?             J@        ������������������������       �                      @        ������������������������       �                     I@        B       C                    #@�3Ea�$�?[            @a@        ������������������������       �                     @        D       {                   �R@���>���?W            �`@       E       v                    �?���A���?V            ``@       F       G                    :@ ���$�?S            �_@        ������������������������       �        	             0@        H       I                    �?�MI8d�?J            �[@        ������������������������       �                     �?        J       u                    �?�2����?I            �[@       K       `                 `fF:@.p����?C            @Y@       L       M                 `f�)@,�+�C�?%            �K@        ������������������������       �                     3@        N       _                   �E@�����H�?             B@       O       V                    @@PN��T'�?             ;@        P       U                    1@��S�ۿ?             .@       Q       T                 �|�=@ףp=
�?             $@        R       S                 �|�<@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        W       Z                   @A@      �?	             (@        X       Y                    1@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        [       ^                   �3@؇���X�?             @       \       ]                   @D@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     "@        a       n                   �B@8����?             G@       b       i                   �C@\X��t�?             7@        c       d                 �|�<@r�q��?             (@        ������������������������       �                     @        e       h                 �|�?@�q�q�?             @       f       g                 `fF<@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        j       k                   �H@���!pc�?	             &@        ������������������������       �                     @        l       m                    K@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        o       p                 ��9L@�nkK�?             7@       ������������������������       �        	             2@        q       r                 �|Y>@z�G�z�?             @        ������������������������       �                      @        s       t                 03�M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        w       x                    �?      �?             @        ������������������������       �                     �?        y       z                   �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        }       �                 Ь�#@���ě)�?�            @y@       ~       �                    �?��!pc�?�            �p@              �                    �?�MI8d�?�            0p@        �       �                 �|�<@H�z�G�?             D@       �       �                    �?�G��l��?             5@       �       �                   �@X�<ݚ�?             2@       �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                 ���@؇���X�?             @        ������������������������       �                     @        �       �                    4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    9@      �?              @        ������������������������       �                     @        �       �                    ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�����?             3@       �       �                 ���@$�q-�?	             *@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 �|Y>@r�q��?             @        ������������������������       �                     @        �       �                    C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �?$@X�M|H�?�            `k@        �       �                 ���@(L���?7            �U@        ������������������������       �                     :@        �       �                 �|Y=@z�G�z�?&             N@        �       �                   �3@���Q��?             4@        ������������������������       �                     @        �       �                    �?      �?	             0@       �       �                    �?��S���?             .@        �       �                 ���@r�q��?             @        ������������������������       �                     @        �       �                   @8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    ;@�q�q�?             "@       �       �                 ���@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?ףp=
�?             D@        �       �                 �|�=@�X�<ݺ?
             2@       �       �                 ���@$�q-�?             *@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 X�,D@��2(&�?             6@       �       �                    �?@�0�!��?             1@       �       �                 �Y�@     ��?             0@        ������������������������       �                     @        �       �                    �?�q�q�?             "@       ������������������������       �����X�?             @        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@�}�+r��?N            �`@        �       �                    �?`���i��?             F@        �       �                 �|Y=@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     A@        �       �                    �?���M�?1            @V@       �       �                   �0@Du9iH��?0            �U@        ������������������������       ��q�q�?             @        �       �                   �;@ ,U,?��?.            �T@        �       �                 @3�!@�����H�?             ;@       �       �                   �:@�LQ�1	�?             7@       �       �                   �2@���N8�?             5@        �       �                 ��Y @؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             ,@        ������������������������       �                      @        ������������������������       �                     @        �       �                 @3�@h�����?             L@        �       �                   �A@ףp=
�?             $@        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                 �|Y?@��<b�ƥ?             G@       �       �                 �|Y=@�nkK�?             7@        ������������������������       �                     @        �       �                 ��) @�IєX�?
             1@       ������������������������       �                     (@        �       �                 pf� @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        ������������������������       �                     @        �       �                   �1@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �                          �?��X��?[            �a@        �       	                   �?� ���?,            @P@       �       �                 @�+@�&!��?            �E@        �       �                    �?ףp=
�?             $@       �       �                 ��&@�����H�?             "@        �       �                 �[$@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�'�=z��?            �@@        ������������������������       �                      @        �       �                    �?`՟�G��?             ?@        �       �                    �?z�G�z�?	             .@       �       �                    �?�q�q�?             "@       �       �                  S�2@      �?             @       �       �                   �-@���Q��?             @        ������������������������       �                      @        �       �                 �|Y6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �                          �?     ��?             0@       �                       03�1@���Q��?             $@       �                           @�q�q�?             @       �       �                 ���.@      �?             @        ������������������������       �                     �?                               �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                              @3�2@r�q��?             @                              ��/@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        
                      `f�8@��2(&�?             6@                                �/@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@              "                   @DE��2{�?/            �R@                             �T)D@`�Q��?"             I@                                �?>��C��?            �E@        ������������������������       �                     @                              ���*@�?�'�@�?             C@                                 )@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                 #@�C��2(�?            �@@        ������������������������       �                      @                                 �?�g�y��?             ?@       ������������������������       �                     ;@                                 �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                 ;@؇���X�?             @        ������������������������       �                     @               !                   >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     9@        �*       h�h))��}�(h,h/h0M#KK��h2h3h4hVh<�h=Kub������������Q�Ȟ���?^-n����?T��_:�?Vx���?L�Ϻ��?�Y7�"��?              �?XG��).�?T\2�h�?�������?�������?�Q����?
ףp=
�?�������?ZZZZZZ�?���Q��?R���Q�?t�E]t�?��.���?UUUUUU�?�������?              �?۶m۶m�?�$I�$I�?              �?333333�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?                      �?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?333333�?�������?              �?      �?              �?      �?      �?                      �?      �?        �������?�������?      �?              �?      �?              �?      �?        ���6��?�� ���?(�����?�k(���?�}A_��?���/��?a���{�?��=���?^Cy�5�?(������?              �?�؉�؉�?ى�؉��?      �?        F]t�E�?]t�E�?      �?      �?              �?      �?                      �?              �?�m۶m��?%I�$I��?      �?      �?      �?      �?      �?                      �?      �?                      �?;�;��?O��N���?      �?                      �?����7��?��,d!�?              �?O�;���?�RKE,�?�eDP�?�i��?�n���v�?�D"�H$�?      �?        ��L���?L�Ϻ��?      �?        ��7�}��?� O	��?�2|#
L�?:5r���?�}��7��?��)A��?      �?        �q�q�?�q�q�?&���^B�?h/�����?�������?�?�������?�������?      �?      �?      �?                      �?      �?              �?              �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?        d!Y�B�?8��Moz�?��Moz��?!Y�B�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?              �?F]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?              �?      �?        �Mozӛ�?d!Y�B�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?^?[���?��N̓�?�.�袋�?�E]t��?��L���?L�Ϻ��?333333�?ffffff�?1�0��?��y��y�?�q�q�?r�q��?�������?�������?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?              �?      �?              �?      �?              �?        ^Cy�5�?Q^Cy��?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?UUUUUU�?      �?              �?      �?              �?      �?        ��QNG9�?\cq��5�?⎸#��?w�qG��?      �?        �������?�������?333333�?�������?      �?              �?      �?�������?�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?                      �?      �?        �������?�������?��8��8�?�q�q�?�؉�؉�?;�;��?      �?              �?      �?      �?        ��.���?t�E]t�?ZZZZZZ�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?      �?      �?      �?              �?        �5��P�?(�����?F]t�E�?F]t�E�?�������?�������?              �?      �?              �?        ��^����?�E(B�?qG�w��?w�qGܱ?UUUUUU�?UUUUUU�?��ˊ��?��FS�׮?�q�q�?�q�q�?��Moz��?Y�B��?��y��y�?�a�a�?۶m۶m�?�$I�$I�?              �?      �?              �?                      �?      �?        �m۶m��?�$I�$I�?�������?�������?      �?        UUUUUU�?UUUUUU�?��7��M�?d!Y�B�?�Mozӛ�?d!Y�B�?      �?        �?�?      �?        �������?�������?              �?      �?              �?              �?        �������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        n۶m۶�?%I�$I��?�����?�ȍ�ȍ�?S֔5eM�?֔5eMY�?�������?�������?�q�q�?�q�q�?      �?      �?              �?      �?                      �?              �?|���?|��|�?      �?        �s�9��?�1�c��?�������?�������?UUUUUU�?UUUUUU�?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��.���?t�E]t�?      �?      �?      �?                      �?      �?        ,�Œ_,�?O贁N�?��(\���?{�G�z�?$�;��?qG�w��?              �?������?y�5���?333333�?�������?              �?      �?        ]t�E�?F]t�E�?              �?��{���?�B!��?      �?              �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ThG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       j                     @<C�`��?�           8�@                                   �?�/DK)��?�            t@                                   �?����=O�?R             b@                                 �6@�IєX�?4            �Y@                                   �?�+$�jP�?             ;@                                 �J@�J�4�?             9@              
                   �9@      �?             8@               	                   �4@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                  @B@P���Q�?             4@       ������������������������       �                     0@                                  �'@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                ��m1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �H@�}��L�?$            �R@       ������������������������       �                     Q@                                83F@؇���X�?             @                                ���;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �E@                                   %@�GN�z�?s             f@        ������������������������       �                     @               5                    �?4>���?n             e@               *                  �>@�Gi����?            �B@                #                   �;@�r����?             .@        !       "                     �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        $       %                   �@@$�q-�?	             *@        ������������������������       �                     @        &       )                     �?؇���X�?             @       '       (                    <@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        +       4                    I@8�A�0��?             6@       ,       -                   �4@������?             1@        ������������������������       �                      @        .       3                    �?�r����?             .@       /       2                 `��I@      �?              @        0       1                 `f�A@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        6       U                     �?��2(&�?R            �`@        7       8                    �?��<b���?)            @Q@        ������������������������       �                      @        9       T                    �?��ga�=�?(            �P@       :       ;                   �<@z�G�z�?'            @P@        ������������������������       �                     @        <       O                   �G@f>�cQ�?%            �N@       =       >                 �|Y>@�ʈD��?            �E@        ������������������������       �        
             .@        ?       H                    �?؇���X�?             <@       @       G                   �F@ףp=
�?             4@       A       B                 �̌/@z�G�z�?             $@        ������������������������       �                     @        C       D                   @@@���Q��?             @        ������������������������       �                      @        E       F                   �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     $@        I       J                 `f�K@      �?              @        ������������������������       �                     @        K       L                 03�M@�q�q�?             @        ������������������������       �                     �?        M       N                    E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        P       S                  i?@�E��ӭ�?
             2@        Q       R                    K@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @        V       i                    �?���N8�?)            �O@       W       X                    �?=QcG��?             �G@        ������������������������       �                      @        Y       h                   �*@��S�ۿ?            �F@       Z       g                    G@�C��2(�?            �@@       [       `                 `fF)@ �Cc}�?             <@       \       _                   �7@�X�<ݺ?             2@        ]       ^                    &@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             *@        a       f                    B@z�G�z�?             $@       b       c                 �|�<@�����H�?             "@       ������������������������       �                     @        d       e                 �|�=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �        	             0@        k       �                 03�7@x�����?�            `x@       l       �                    �?$6HZl�?�            @u@        m       x                 �̌@8�A�0��?/            �P@        n       w                    @      �?             8@       o       p                    8@�����?             3@        ������������������������       �                     @        q       v                    �?      �?
             (@       r       u                    �?      �?              @       s       t                 ���@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        y       �                 �|�<@      �?             E@       z                           �?���|���?             6@        {       |                    �?z�G�z�?             @        ������������������������       �                      @        }       ~                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �*@������?             1@       �       �                 ��&@���|���?	             &@       �       �                    �?�<ݚ�?             "@       �       �                    �?      �?              @        �       �                 �̼!@      �?             @        ������������������������       �                      @        �       �                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��Q��?             4@        �       �                    �?����X�?             @       �       �                 P�h2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��� @8�Z$���?
             *@        ������������������������       �                     �?        �       �                   �>@�8��8��?	             (@       ������������������������       �                      @        �       �                    �?      �?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                 ���0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?����l��?�             q@       �       �                 �?�@P��4���?�            �o@       �       �                 �Y�@�L#���?P            �`@        �       �                    �?      �?             H@        �       �                 ��y@8�Z$���?             :@        ������������������������       �                     @        �       �                 ���@"pc�
�?             6@        �       �                   �7@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        �       �                   �5@�<ݚ�?             "@        ������������������������       �                     �?        �       �                 �|=@      �?              @        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                 ���@�C��2(�?             6@       ������������������������       �                     4@        ������������������������       �                      @        �       �                    �? qP��B�?5            �U@       �       �                 ��]@�Ń��̧?3             U@       ������������������������       �                    �H@        �       �                 �Yu@ >�֕�?            �A@        �       �                    >@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     >@        ������������������������       �                      @        �       �                    �?����\�?M            @^@       �       �                 ��q1@r�q��??             X@       �       �                   `!@*
;&���?<             W@       �       �                    �?d��0u��?(             N@        ������������������������       �                     �?        �       �                   �3@��$�4��?'            �M@        �       �                 0S5 @      �?             (@       �       �                    1@���Q��?             $@        ������������������������       ����Q��?             @        �       �                   �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        �       �                 @3�@��0{9�?!            �G@        �       �                    :@      �?              @        ������������������������       �                     @        �       �                   �?@���Q��?             @        ������������������������       �                     �?        �       �                   �A@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                 �|Y<@��-�=��?            �C@        �       �                   �:@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        �       �                 ��) @h�����?             <@       ������������������������       �                     4@        �       �                 ��y @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �<@      �?             @@       ������������������������       �                     3@        �       �                 �|Y=@$�q-�?	             *@        �       �                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?      �?             @       �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��Y)@z�G�z�?             9@        �       �                    8@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�}�+r��?             3@       ������������������������       �                     ,@        �       �                  �v6@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|Y?@�\��N��?             3@       �       �                 ��\"@�	j*D�?             *@        ������������������������       �                      @        �       �                    �?"pc�
�?             &@        ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                    $@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �                           ?@ "��u�?             I@       �       �                     @ ���J��?            �C@        �       �                    �?؇���X�?             @       �       �                 �|�3@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @@                                 �?"pc�
�?             &@                                �A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                              ��A>@؇���X�?             @        ������������������������       �                     @                                 @      �?             @        ������������������������       �                      @        	      
                  �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������܍�W�?/�F�JP�?^
3�O�?��z���?��RA�/�?U��K��?�?�?B{	�%��?/�����?{�G�z�?�z�G��?      �?      �?      �?      �?              �?      �?        �������?ffffff�?              �?      �?      �?              �?      �?              �?              �?      �?              �?      �?        O贁N�?�_,�Œ�?              �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?�袋.��?]t�E�?              �?��]�`��?�T�6|��?o0E>��?#�u�)��?�������?�?      �?      �?              �?      �?        �؉�؉�?;�;��?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?              �?      �?              �?        /�袋.�?颋.���?�?xxxxxx�?      �?        �?�������?      �?      �?      �?      �?              �?      �?                      �?              �?      �?        ��.���?t�E]t�?��,d!�?��Moz��?      �?        ��[���?�1���?�������?�������?              �?��!XG�?�u�y���?A_���?�}A_з?      �?        ۶m۶m�?�$I�$I�?�������?�������?�������?�������?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �q�q�?r�q��?      �?      �?              �?      �?              �?                      �?��y��y�?�a�a�?x6�;��?AL� &W�?      �?        �������?�?]t�E�?F]t�E�?%I�$I��?۶m۶m�?��8��8�?�q�q�?�������?�������?              �?      �?              �?        �������?�������?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?              �?        ��o��o�?�A�A�?�������?�������?/�袋.�?颋.���?      �?      �?^Cy�5�?Q^Cy��?              �?      �?      �?      �?      �?�$I�$I�?۶m۶m�?      �?                      �?      �?              �?                      �?      �?      �?]t�E]�?F]t�E�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?xxxxxx�?�?]t�E]�?F]t�E�?9��8���?�q�q�?      �?      �?      �?      �?      �?              �?      �?              �?      �?              �?                      �?              �?      �?        ffffff�?�������?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        ;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?)��?�[�w��?\\\\\\�?�?��@���?g��1��?      �?      �?;�;��?;�;��?      �?        /�袋.�?F]t�E�?;�;��?;�;��?              �?      �?        9��8���?�q�q�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?]t�E�?F]t�E�?      �?                      �?��}A�?�}A_З?��<��<�?�a�a�?      �?        ��+��+�?�A�A�?333333�?�������?      �?                      �?      �?              �?        �T�x?r�?}��7�?�������?UUUUUU�?���,d!�?8��Moz�?�?�������?      �?        #h8����?u_[4�?      �?      �?�������?333333�?333333�?�������?�������?�������?              �?      �?      �?      �?        m�w6�;�?L� &W�?      �?      �?      �?        �������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?}˷|˷�?�A�A�?F]t�E�?t�E]t�?      �?                      �?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?              �?      �?      �?        �؉�؉�?;�;��?      �?      �?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?        �5��P�?(�����?      �?        �������?�������?      �?                      �?y�5���?�5��P�?;�;��?vb'vb'�?      �?        F]t�E�?/�袋.�?              �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �G�z�?���Q��?��-��-�?�A�A�?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?              �?      �?              �?              �?        /�袋.�?F]t�E�?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?      �?              �?      �?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ5�R/hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       ^                    �?t�C�#��?�           8�@               )                     @�T����?�            0p@                                  �? sAr�=�?X            �b@        ������������������������       �                     F@               (                    �?ܾ�z�<�?=             Z@              %                    L@��8��)�?8            �W@                                  6@������?5            @V@                                  @4@r�q��?             >@       	                           :@$�q-�?             :@        
                           �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�nkK�?             7@                                 �*@���N8�?             5@                               `f�)@��S�ۿ?
             .@        ������������������������       �                     @                                  �B@ףp=
�?             $@       ������������������������       �                      @                                   D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                    �?���#�İ?#            �M@                                 �E@ pƵHP�?             J@       ������������������������       �                     F@                                  @F@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        !       $                     �?؇���X�?             @        "       #                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        &       '                   �L@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        *       A                    �?P7Z�U��?C            �[@        +       4                    �?�+e�X�?              I@        ,       -                    �?�>����?             ;@        ������������������������       �                     "@        .       3                    @�����H�?             2@       /       0                 �|�9@�IєX�?
             1@        ������������������������       �                     @        1       2                 ���@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        5       @                   �;@\X��t�?             7@       6       ?                    �?�E��ӭ�?             2@       7       8                    5@      �?             $@        ������������������������       �                      @        9       >                 03�!@      �?              @       :       ;                    8@r�q��?             @       ������������������������       �                     @        <       =                 pff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        B       Y                    �?�'N��?#            �N@       C       N                    �?     ��?             @@       D       E                 @%@��.k���?             1@        ������������������������       �                     @        F       I                 �|�;@�n_Y�K�?	             *@        G       H                    0@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        J       K                 �|Y>@�<ݚ�?             "@        ������������������������       �                     @        L       M                 03�1@      �?             @       ������������������������       �                      @        ������������������������       �                      @        O       R                    �?��S���?
             .@        P       Q                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        S       X                     @      �?             (@       T       U                    0@�q�q�?             "@        ������������������������       �                     @        V       W                    >@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        Z       [                 X��@@ 	��p�?             =@       ������������������������       �                     4@        \       ]                   @C@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        _       r                 �?�@�6�F8)�?#           @|@        `       g                    �?`Ql�R�?W            �a@        a       f                    �?�X�<ݺ?             2@       b       e                 �|Y=@�IєX�?             1@        c       d                   �<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             (@        ������������������������       �                     �?        h       i                 ��@�-.�1a�?I            �^@       ������������������������       �        (            �O@        j       k                    �?(;L]n�?!             N@        ������������������������       �                      @        l       m                 �|Y=@XB���?              M@       ������������������������       �                    �B@        n       q                 �|�=@�����?             5@       o       p                  sW@؇���X�?	             ,@        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     @        s       �                    @z��!���?�            ps@       t       �                 @�:x@BSf���?�            r@       u       v                    ,@��G�<�?�            �q@        ������������������������       �                     ,@        w       �                    @"�m詹�?�            �p@       x       �                     �?� �(���?�            �p@        y       �                    �?�P�����?>             U@       z       �                    �?P��MO�?=            �T@        {       �                    �?¦	^_�?             ?@       |       �                   @H@������?             >@       }       �                   @C@�ՙ/�?             5@       ~       �                 �|Y<@�����?             3@              �                    �?�eP*L��?             &@       �       �                   �7@      �?              @        ������������������������       �                      @        �       �                    �?r�q��?             @       �       �                   �9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �U�X@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?              @       �       �                   @@@r�q��?             @       ������������������������       �                     @        �       �                   �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?���3�E�?'             J@       �       �                   �<@     ��?$             H@        �       �                    7@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @       �       �                 `f�D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���?            �D@       �       �                  i?@������?             >@       �       �                   @>@X�<ݚ�?             2@       �       �                    R@      �?             0@       �       �                    J@����X�?             ,@       �       �                 �|�?@      �?              @        ������������������������       �                     @        �       �                    D@z�G�z�?             @        ������������������������       �                      @        �       �                   @G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        �       �                 `�iJ@"pc�
�?             &@        ������������������������       �                     �?        �       �                   �D@ףp=
�?             $@        �       �                   �B@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?������?r             g@        �       �                    �?���|���?             &@        �       �                 ���/@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 03�-@      �?              @        ������������������������       �                     @        �       �                 �|Y>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     @���(`�?k            �e@        �       �                   �@@Hn�.P��?)             O@       ������������������������       �                     B@        �       �                    �?ȵHPS!�?             :@       �       �                    �?�S����?             3@        ������������������������       �                     �?        �       �                    �?r�q��?             2@       �       �                    ,@z�G�z�?
             .@       �       �                 `f�)@�q�q�?             "@        ������������������������       �                     @        �       �                   �A@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�X�C�?B             \@        ������������������������       �                     @        �       �                 �|Y=@�u��R�??            �Z@       �       �                 0S5 @��x_F-�?             �I@        �       �                 @3�@�q�q�?	             .@        ������������������������       �                     �?        �       �                   �3@X�Cc�?             ,@        �       �                   �1@r�q��?             @       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?4?,R��?             B@       �       �                   �8@r�q��?             >@       ������������������������       �                     4@        �       �                   �;@      �?             $@        ������������������������       �                     @        �       �                   �<@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�h����?             L@       �       �                   �>@��<D�m�?            �H@       ������������������������       �                     7@        �       �                   �?@ȵHPS!�?             :@        ������������������������       �                     �?        �       �                   �@@HP�s��?             9@        ������������������������       ��q�q�?             @        �       �                 @3�@���7�?	             6@        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @���7�?             6@        �       �                    @؇���X�?             @        ������������������������       �                      @        �       �                    @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub���������������td�@�?��7a~�?� U���?�ո��?*�Y7�"�?�`�|��?              �?vb'vb'�?�;�;�?br1���?�Q�٨��?B�P�"�?ؽ�u�{�?UUUUUU�?�������?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?      �?                      �?d!Y�B�?�Mozӛ�?�a�a�?��y��y�?�?�������?              �?�������?�������?              �?      �?      �?      �?                      �?              �?              �?      �?      �?              �?      �?        'u_[�?��N��?;�;��?'vb'vb�?              �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?�������?333333�?      �?                      �?              �?Nq��$�?c��2��?���Q��?R���Q�?h/�����?�Kh/��?              �?�q�q�?�q�q�?�?�?              �?;�;��?�؉�؉�?      �?                      �?      �?        ��Moz��?!Y�B�?r�q��?�q�q�?      �?      �?      �?              �?      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?                      �?      �?        �����?ާ�d��?      �?      �?�������?�?      �?        ى�؉��?;�;��?      �?      �?              �?      �?        �q�q�?9��8���?              �?      �?      �?              �?      �?        �?�������?UUUUUU�?UUUUUU�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        ������?�{a���?      �?        9��8���?�q�q�?              �?      �?        04��A�?B�/4��?}g���Q�?W�+�ɕ?��8��8�?�q�q�?�?�?�������?�������?      �?                      �?      �?              �?        {����z�?�h
���?      �?        �������?�?      �?        GX�i���?�{a���?      �?        =��<���?�a�a�?۶m۶m�?�$I�$I�?              �?      �?              �?        m�%�/j�?J�hAW�?躍`3�?`�}2��?�m�`�?��I��?              �?ZO�m���?�®I.A�?�f�P���?�dn��i�?��y��y�?�0�0�?��7�:��?���ˊ��?��Zk���?�RJ)���?wwwwww�?�?�<��<��?�a�a�?Q^Cy��?^Cy�5�?t�E]t�?]t�E�?      �?      �?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?      �?                      �?O��N���?b'vb'v�?      �?      �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?�������?�������?              �?      �?                      �?28��1�?8��18�?wwwwww�?�?r�q��?�q�q�?      �?      �?�m۶m��?�$I�$I�?      �?      �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?      �?        /�袋.�?F]t�E�?              �?�������?�������?      �?      �?      �?                      �?      �?              �?                      �?��g�`��?к����?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?              �?      �?              �?      �?        g��o��?Ȥx�L��?t�9�s�?�c�1ƨ?      �?        ��N��N�?�؉�؉�?(������?^Cy�5�?      �?        �������?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?              �?        �$I�$I�?n۶m۶�?      �?        �@�Ե�?7��XQ�?�������?�?UUUUUU�?UUUUUU�?      �?        %I�$I��?�m۶m��?UUUUUU�?�������?      �?      �?              �?      �?        �8��8��?r�q��?�������?UUUUUU�?      �?              �?      �?              �?�m۶m��?�$I�$I�?      �?                      �?      �?        �$I�$I�?۶m۶m�?��S�r
�?և���X�?      �?        ��N��N�?�؉�؉�?              �?q=
ףp�?{�G�z�?UUUUUU�?UUUUUU�?�.�袋�?F]t�E�?              �?      �?              �?              �?                      �?�.�袋�?F]t�E�?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�%hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM)hjh))��}�(h,h/h0M)��h2h3h4hph<�h=Kub������       d                    �?>AU`�z�?�           8�@               %                    �?xh&���?z             h@                                ���@�����H�?5            @T@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�:�^���?3            �S@              	                    �?@3����?"             K@       ������������������������       �                     ?@        
                         S�-@�nkK�?             7@                                    @r�q��?             @        ������������������������       �                      @                                �|Y6@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     1@               $                    �?      �?             8@              !                    E@��<b���?             7@                                   @�S����?             3@        ������������������������       �                     @                                    @      �?             (@                                  �?�z�G��?             $@                                  �?      �?              @                                  �?�q�q�?             @        ������������������������       �                     �?                                �|Y3@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        "       #                      @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        &       '                    �?����X��?E             \@        ������������������������       �                     @        (       Q                 ���=@�G�.o�?C            @[@       )       D                    �?b:�&���?3            �T@       *       1                   �6@�D��?            �H@        +       0                    �?����X�?             @       ,       -                    '@�q�q�?             @        ������������������������       �                     �?        .       /                 ��y@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        2       C                 м;4@��s����?             E@       3       B                 �|Y?@������?             >@       4       5                   �8@���|���?             6@        ������������������������       �                     @        6       A                 03�-@D�n�3�?             3@       7       @                    �?d}h���?             ,@       8       9                 ���@      �?	             (@        ������������������������       �                     @        :       =                   @@և���X�?             @       ;       <                 �|=@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        >       ?                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        E       N                    �?�IєX�?             A@       F       M                 ��(@h�����?             <@       G       L                 X��A@�X�<ݺ?             2@       H       K                    �?��S�ۿ?	             .@       I       J                 ���@�8��8��?             (@        ������������������������       �                     @        ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        O       P                 �|�2@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        R       ]                 @��V@      �?             :@       S       \                 ��UO@����X�?	             ,@       T       [                    �?X�<ݚ�?             "@       U       Z                   @J@����X�?             @       V       W                    �?r�q��?             @        ������������������������       �                     @        X       Y                     �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ^       c                    �?      �?             (@       _       `                 X�,@@      �?              @        ������������������������       �                     @        a       b                   @E@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        e       (                   @~�hP��?O           0�@       f                          �?b�^y,�?A            @       g       �                 �|�=@:�{0��?�            �w@       h       s                     �?�5��
J�?�            �l@        i       j                   @>@�LQ�1	�?             7@        ������������������������       �                     @        k       l                    �?���y4F�?
             3@        ������������������������       �                      @        m       n                   �D@���|���?             &@        ������������������������       �                     @        o       p                    �?և���X�?             @        ������������������������       �                      @        q       r                    7@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        t       �                     @@w�h��?�            �i@        u       z                    �?��i#[�?             E@        v       w                    1@$�q-�?
             *@       ������������������������       �                      @        x       y                   �7@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        {       �                    &@XB���?             =@        |       }                    @ףp=
�?             $@        ������������������������       �                     @        ~                           5@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        �       �                    �?�2����?g            �d@        �       �                 ���@`՟�G��?             ?@        ������������������������       �                     @        �       �                  �#@�q�q�?             8@       �       �                   �3@$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        �       �                 �|�;@�eP*L��?             &@       �       �                 @�)@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �T)D@p^H�&m�?T            �`@       �       �                    �?,mG����?Q             `@       �       �                 �?�@4Jı@�?O            �_@        �       �                 �?$@���#�İ?&            �M@       �       �                 ��@ 	��p�?             =@       �       �                    7@ �q�q�?             8@       ������������������������       �        	             *@        �       �                   �8@�C��2(�?             &@        �       �                 `fF@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 �|Y8@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     >@        �       �                    �?�G�V�e�?)             Q@       �       �                 @3�!@�?�<��?&            @P@       �       �                 �|Y<@��s����?             E@       �       �                   �:@      �?             <@       �       �                 0S5 @�J�4�?             9@       �       �                 @3�@������?
             1@        ������������������������       �                     @        �       �                   �4@���|���?             &@       �       �                    1@և���X�?             @        ������������������������       �                      @        �       �                   �2@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��) @@4և���?
             ,@       ������������������������       �                     (@        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        �       �                 �|�8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    ;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �K@���=A�?k             c@       �       �                    �?���|���?]            �`@        �       �                    �?z�G�z�?             D@       �       �                   @B@؇���X�?             5@        ������������������������       �                     &@        �       �                   �C@�z�G��?	             $@        ������������������������       �                      @        �       �                   @"@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @@�d�����?             3@        ������������������������       �                     @        �       �                     �?      �?
             0@        ������������������������       �                     @        �       �                     @�<ݚ�?             "@        �       �                   �E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��Y.@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �G@�㙢�c�?A             W@       �       �                 0�K@�o��gn�?<            �T@       �       �                   �?@�C��2(�?7            @S@        �       �                    �?�θ�?	             *@       �       �                   �>@      �?             (@       �       �                     @      �?              @        ������������������������       �                     @        �       �                 �̌!@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                      @      �?             @        ������������������������       �                     �?        �       �                 pff@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��$:@      �?.             P@       �       �                   @@@@3����?&             K@        �       �                    �?      �?              @       �       �                   �@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      G@        �       �                   @C@�z�G��?             $@        ������������������������       �                      @        �       �                 `f�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �D@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �H@X�<ݚ�?             "@        ������������������������       �                      @        �       �                    3@և���X�?             @        ������������������������       �                      @        �       �                 03�D@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �                          @S@ףp=
�?             4@       �       �                     �?�}�+r��?             3@       �       �                 `vo=@�8��8��?             (@       �       �                   �M@�����H�?             "@        �       �                   �L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?              %                   @>n�T��?E             ]@                                �?�VbbP�??            �Z@                                �?D|U��@�?%            �P@        ������������������������       �                     >@              	                    @����>�?            �B@                                @�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        
                         @X�Cc�?
             ,@        ������������������������       �                     @                                 A@ףp=
�?             $@       ������������������������       �                     @                                �E@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                              `ff.@�z�G��?             D@        ������������������������       �                      @              $                   �?      �?             @@             #                03c@�q�q�?             >@             "                   @�q�q�?             8@             !                `��S@�eP*L��?             6@                                 :@�q�q�?             2@                                0@��
ц��?
             *@        ������������������������       �                     �?                                  @�q�q�?	             (@                                �3@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                 +@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        &      '                     @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     4@        �*       h�h))��}�(h,h/h0M)KK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?b6�5��?�d�x��?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?        �o��o��?� � �?h/�����?���Kh�?              �?d!Y�B�?�Mozӛ�?UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?      �?      �?��Moz��?��,d!�?^Cy�5�?(������?              �?      �?      �?333333�?ffffff�?      �?      �?UUUUUU�?UUUUUU�?              �?�������?333333�?      �?                      �?      �?      �?              �?      �?                      �?              �?      �?      �?              �?      �?              �?        I�$I�$�?n۶m۶�?              �?z|���?��p�?�b��7�?o4u~�!�?������??4և���?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?                      �?              �?z��y���?�a�a�?wwwwww�?�?]t�E]�?F]t�E�?      �?        l(�����?(������?I�$I�$�?۶m۶m�?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?              �?        �?�?�m۶m��?�$I�$I�?��8��8�?�q�q�?�������?�?UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?      �?              �?              �?        �������?UUUUUU�?      �?                      �?      �?      �?�$I�$I�?�m۶m��?�q�q�?r�q��?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?      �?      �?      �?      �?      �?        �������?333333�?              �?      �?              �?        S�n0�?�Y7�"��?����H��?�dn}�?C�E4�?��y�t��?�,d!Y�?�Mozӛ�?d!Y�B�?Nozӛ��?      �?        (������?6��P^C�?              �?F]t�E�?]t�E]�?              �?�$I�$I�?۶m۶m�?      �?        �������?333333�?      �?                      �?HZ�<��?ᖚ���?�a�a�?�<��<��?;�;��?�؉�؉�?              �?�������?�������?      �?                      �?GX�i���?�{a���?�������?�������?      �?        �������?UUUUUU�?              �?      �?              �?        ��7�}��?� O	��?�1�c��?�s�9��?              �?�������?�������?�؉�؉�?;�;��?              �?      �?        ]t�E�?t�E]t�?�������?UUUUUU�?              �?      �?                      �?`���@��?��[�ո?QW�uE�?uE]QWԵ?O���t:�?��b�X,�?��N��?'u_[�?������?�{a���?�������?UUUUUU�?      �?        ]t�E�?F]t�E�?      �?      �?              �?      �?              �?        �������?�������?      �?              �?      �?      �?        �������?�������?�����? �����?z��y���?�a�a�?      �?      �?�z�G��?{�G�z�?xxxxxx�?�?      �?        ]t�E]�?F]t�E�?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?      �?      �?              �?                      �?n۶m۶�?�$I�$I�?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?        333333�?�������?              �?      �?        ��P^Cy�?�P^Cy�?]t�E]�?F]t�E�?�������?�������?�$I�$I�?۶m۶m�?              �?333333�?ffffff�?      �?              �?      �?      �?                      �?y�5���?Cy�5��?      �?              �?      �?              �?�q�q�?9��8���?      �?      �?              �?      �?        �������?�������?      �?                      �?�7��Mo�?d!Y�B�?rY1P��?�7�:���?]t�E�?F]t�E�?ى�؉��?�؉�؉�?      �?      �?      �?      �?      �?        �������?�������?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?���Kh�?h/�����?      �?      �?۶m۶m�?�$I�$I�?              �?      �?              �?              �?        ffffff�?333333�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �q�q�?r�q��?              �?�$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?        �������?�������?�5��P�?(�����?UUUUUU�?UUUUUU�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?                      �?��{a�?,�4�rO�?�#蝺�?n����?�rv��?Xc"=P9�?              �?���L�?�u�)�Y�?d!Y�B�?�Mozӛ�?      �?                      �?%I�$I��?�m۶m��?              �?�������?�������?      �?              �?      �?              �?      �?        ffffff�?333333�?      �?              �?      �?UUUUUU�?UUUUUU�?�������?�������?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?�;�;�?�؉�؉�?              �?�������?�������?�������?333333�?              �?      �?        �m۶m��?�$I�$I�?              �?      �?              �?                      �?      �?              �?                      �?�q�q�?�q�q�?              �?      �?              �?        �       ubhhubehhub.