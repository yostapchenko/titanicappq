��]      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�_sklearn_version��1.5.1�ub�n_estimators�Kd�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK*�verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hNhG        �feature_names_in_��joblib.numpy_pickle��NumpyArrayWrapper���)��}�(�subclass��numpy��ndarray����shape�K���order��C��dtype�h-�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�
allow_mmap���numpy_array_alignment_bytes�Kub�cnumpy.core.multiarray
_reconstruct
q cnumpy
ndarray
qK �qc_codecs
encode
qX   bqX   latin1q�qRq�qRq	(KK�q
cnumpy
dtype
qX   O8q���qRq(KX   |qNNNJ����J����K?tqb�]q(X   PclassqX   SexqX   AgeqX   ParchqX   FareqX   Embarkedqetqb.��       �n_features_in_�K�
_n_samples�M��
n_outputs_�K�classes_�h))��}�(h,h/h0K��h2h3h4h6�i8�����R�(K�<�NNNJ����J����K t�bh<�h=Kub�               ��       �
n_classes_�K�_n_samples_bootstrap�M��
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJf��_hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4h6�f8�����R�(KhHNNNJ����J����K t�bh<�h=Kub��������������              �?��       hJ�numpy.core.multiarray��scalar���hGC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub���       �k      K��R�}�(hK�
node_count�M�nodes�h))��}�(h,h/h0M��h2h3h4h6�V64�����R�(Kh:N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(hqh6�i8�����R�(KhHNNNJ����J����K t�bK ��hrh}K��hsh}K��hthVK��huhVK ��hvh}K(��hwhVK0��hxh6�u1�����R�(Kh:NNNJ����J����K t�bK8��uK@KKt�bh<�h=Kub���       R                    �?���*1�?�           8�@                                    @�U>�� �?�             o@                                 �&@ȥ�fzR�?Y             a@                                  �J@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @                                   @X�GP>��?S            �_@        ������������������������       �                      @        	       
                   �B@`2U0*��?R            @_@       ������������������������       �        :            @V@                                �QD@4?,R��?             B@                                   �?�n_Y�K�?	             *@                                  �?�q�q�?             (@        ������������������������       �                      @                                 ��9@�z�G��?             $@                                   �?      �?              @        ������������������������       �                      @                                  �,@r�q��?             @                                   D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@               -                    �?��7Y��?G            �[@               $                    �?H�V�e��?             A@                                 �-@�>����?             ;@                                �&�)@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                #                 ���@���7�?             6@        !       "                 �Y�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@        %       ,                    @����X�?             @       &       +                    �?�q�q�?             @       '       (                    '@      �?             @        ������������������������       �                     �?        )       *                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        .       I                    �?:���u��?/            @S@       /       <                 ��&@θ	j*�?              J@       0       5                   �3@@�0�!��?             A@        1       4                 �&B@r�q��?             @        2       3                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        6       7                   �9@h�����?             <@       ������������������������       �                     ,@        8       ;                 @3�@@4և���?             ,@        9       :                 �?�@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        =       >                    '@b�2�tk�?             2@        ������������������������       �                     @        ?       @                   �6@      �?
             ,@        ������������������������       �                     @        A       F                    �?�z�G��?             $@       B       C                 �|Y>@؇���X�?             @        ������������������������       �                     @        D       E                    @@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        G       H                   �;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        J       K                 @34@HP�s��?             9@        ������������������������       �                     �?        L       Q                    @ �q�q�?             8@       M       P                    @      �?	             0@        N       O                 ��T?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                      @        S       �                     �?��V�[�?$           �|@        T       �                    �?�U���?F             _@       U       t                  x#J@Ru߬��?A            �\@       V       W                 �|�<@ٜSu��?(            @Q@        ������������������������       �                     @        X       o                   �D@     ��?%             P@       Y       h                   �@@4�B��?            �B@       Z       a                    �?�㙢�c�?             7@        [       `                 ��2>@r�q��?             @       \       _                 �|�=@�q�q�?             @       ]       ^                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        b       g                 �|Y>@@�0�!��?
             1@       c       d                 `fF<@z�G�z�?             .@        ������������������������       �                     @        e       f                   �>@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        i       l                    �?և���X�?             ,@        j       k                   �A@      �?              @       ������������������������       �                     @        ������������������������       �                     @        m       n                   �B@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        p       s                   @J@�>����?             ;@        q       r                   �G@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �        	             ,@        u       �                   @I@��S���?            �F@       v       �                    �?�n_Y�K�?            �C@       w       x                   �8@�q�q�?             >@        ������������������������       �                     @        y       |                    �?������?             ;@       z       {                   �H@@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        }       �                   �B@��
ц��?             *@        ~                        �|Y>@z�G�z�?             @        ������������������������       �                      @        �       �                 `f�K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �E@      �?              @        ������������������������       �                     @        �       �                   �G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �7@X�<ݚ�?             "@        ������������������������       �                      @        �       �                 �̾w@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �̰f@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                     @����?�            0u@        �       �                   �)@؇���X�?4            �Q@        �       �                    �?`2U0*��?             9@        ������������������������       �                     @        �       �                    4@���N8�?             5@        �       �                   �2@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �        
             0@        �       �                    �?z�G�z�?$            �F@       �       �                   �*@      �?             @@       �       �                 �|�<@������?             1@        ������������������������       �                     @        �       �                 �|�=@���|���?	             &@        ������������������������       �                     �?        �       �                   �F@�z�G��?             $@       �       �                    @@      �?              @        ������������������������       �                     �?        �       �                   �C@և���X�?             @       �       �                   �A@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     .@        �       �                    ,@�n_Y�K�?
             *@        ������������������������       �                     @        ������������������������       �                      @        �       �                 ��-@܉���?�            �p@       �       �                    &@LܤK���?�            �j@        ������������������������       �                      @        �       �                    �?��au���?�            �j@        �       �                 ���@�n`���?             ?@        �       �                 �|�9@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?      �?             4@       �       �                   �5@�E��ӭ�?             2@        ������������������������       �                      @        �       �                 �|�=@     ��?             0@       �       �                 ��� @      �?	             (@       �       �                   @:@�q�q�?             "@        ������������������������       �                     �?        �       �                   @@      �?              @       ������������������������       ��q�q�?             @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?���fu�?q            �f@       �       �                 @3�@��;M��?o            @f@       �       �                    �?�}�+r��?H            �\@        �       �                 �|Y=@�����H�?             ;@        ������������������������       �                     @        ������������������������       �                     8@        �       �                   �7@XB���?;            �U@        ������������������������       �                     A@        �       �                 �|Y>@ �h�7W�?%            �J@       �       �                 �?$@�����H�?             ;@        �       �                 pf�@d}h���?
             ,@       �       �                 ���@�C��2(�?             &@        �       �                   �8@z�G�z�?             @        �       �                 �&b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     :@        �       �                   �3@     ��?'             P@        �       �                   �1@�t����?
             1@        �       �                   �0@�<ݚ�?             "@       �       �                 pFD!@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `�8"@      �?              @       �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                 ��) @dP-���?            �G@        ������������������������       �        	             .@        �       �                 ��y @      �?             @@        ������������������������       �                     �?        �       �                 ���"@��a�n`�?             ?@       �       �                 @3�!@�}�+r��?             3@       �       �                 �|Y<@��S�ۿ?             .@        �       �                   �:@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �       �                 `�X#@r�q��?             (@       �       �                   �<@�<ݚ�?             "@        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �                           0@���!pc�?$            �K@        �       �                    �?�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @                                 �?:	��ʵ�?            �F@                                �2@      �?             @        ������������������������       �                     �?                              м;4@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                              �T�I@�p ��?            �D@                                �?`Jj��?             ?@        	      
                03�6@�r����?             .@       ������������������������       �                     (@                              03�7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@                              �|�>@���Q��?             $@                             �|�;@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �1       �values�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�����`l����??'��d�?[k���Z�?SJ)��R�?T{N���?}�06��?333333�?ffffff�?              �?      �?        ���p8�?����x<�?      �?        {�G�z�?���Q��?              �?r�q��?�8��8��?ى�؉��?;�;��?�������?�������?      �?        333333�?ffffff�?      �?      �?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?                      �?              �?�+c���?\�9	ą�?ZZZZZZ�?iiiiii�?h/�����?�Kh/��?�������?�������?              �?      �?        F]t�E�?�.�袋�?UUUUUU�?UUUUUU�?              �?      �?                      �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        dj`��?qV~B���?�؉�؉�?�N��N��?ZZZZZZ�?�������?UUUUUU�?�������?      �?      �?              �?      �?                      �?�m۶m��?�$I�$I�?      �?        n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        9��8���?�8��8��?              �?      �?      �?      �?        333333�?ffffff�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        q=
ףp�?{�G�z�?              �?�������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        u5`:�?+�+��?c�1��?�9�s��?�>����??���#�?s��\;0�?%~F���?              �?      �?      �?�Y7�"��?L�Ϻ��?�7��Mo�?d!Y�B�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        ZZZZZZ�?�������?�������?�������?      �?              �?      �?              �?      �?              �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?        UUUUUU�?�������?              �?      �?        �Kh/��?h/�����?;�;��?;�;��?      �?                      �?      �?        �������?�?ى�؉��?;�;��?UUUUUU�?UUUUUU�?      �?        {	�%���?B{	�%��?�$I�$I�?n۶m۶�?              �?      �?        �؉�؉�?�;�;�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?r�q��?�q�q�?              �?�m۶m��?�$I�$I�?      �?                      �?      �?        333333�?ffffff�?              �?      �?        "��x�?x�!���?۶m۶m�?�$I�$I�?���Q��?{�G�z�?      �?        ��y��y�?�a�a�?�������?�������?      �?              �?      �?      �?        �������?�������?      �?      �?xxxxxx�?�?      �?        ]t�E]�?F]t�E�?              �?ffffff�?333333�?      �?      �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?              �?        ;�;��?ى�؉��?              �?      �?        ��k�z�?�Q���?�B�(���?蝺���?              �?0��>���?~�	�[�?�9�s��?�c�1��?]t�E�?F]t�E�?              �?      �?              �?      �?�q�q�?r�q��?              �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?              �?        �8x�Y�?g;>)7�?զ6��M�?Y�JV���?�5��P�?(�����?�q�q�?�q�q�?              �?      �?        GX�i���?�{a���?      �?        ��sHM0�?"5�x+��?�q�q�?�q�q�?I�$I�$�?۶m۶m�?]t�E�?F]t�E�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?             ��?      �?�������?�������?9��8���?�q�q�?333333�?�������?              �?      �?              �?              �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        �����F�?W�+�ɵ?      �?              �?      �?              �?�s�9��?�c�1Ƹ?�5��P�?(�����?�������?�?�������?�������?      �?                      �?      �?              �?        �������?UUUUUU�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        F]t�E�?t�E]t�?333333�?ffffff�?      �?                      �?��O��O�?l�l��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        Q��+Q�?��+Q��?���{��?�B!��?�������?�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        333333�?�������?۶m۶m�?�$I�$I�?              �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�=�KhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������                           @\AK"���?�           8�@                                ��*4@���"͏�?            �B@        ������������������������       �        	             0@                                �̌5@և���X�?             5@        ������������������������       �                     @                                  �C@�t����?             1@              
                    �?�C��2(�?             &@               	                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@                                    @�q�q�?             @                               p"$X@      �?             @        ������������������������       �                     �?                                �(\�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @               x                     @H�g����?�           �@               +                    �?� k����?�            s@               *                    �?H�Swe�?Q            @_@                                 �B@���M�?9            @V@                                 �6@��.N"Ҭ?)            @Q@                                ��m1@�C��2(�?             6@       ������������������������       �                     3@                                   ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �G@                                  �C@z�G�z�?             4@        ������������������������       �                     �?                %                     �?�S����?             3@       !       $                   �I@؇���X�?
             ,@        "       #                   �H@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        &       '                   �E@z�G�z�?             @       ������������������������       �                     @        (       )                   �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     B@        ,       o                    �?DG��L�?p            �f@       -       :                 ��$:@��A��?^            �b@        .       /                    �? ��ʻ��?.             Q@        ������������������������       �                     @        0       1                 `f�)@ ������?*            �O@        ������������������������       �                     ?@        2       3                     �?      �?             @@        ������������������������       �                     @        4       9                   �*@XB���?             =@       5       6                   @D@�IєX�?             1@       ������������������������       �                     (@        7       8                   �F@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     (@        ;       P                    �?     ��?0             T@        <       O                    J@�q�����?             9@       =       >                 �ܵ<@���Q��?             4@        ������������������������       �                      @        ?       @                   �8@�q�q�?             2@        ������������������������       �                      @        A       H                 0��G@      �?             0@        B       C                  Y>@      �?             @        ������������������������       �                      @        D       E                  �>@      �?             @        ������������������������       �                      @        F       G                 `f�A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       J                 �|Y<@ףp=
�?             $@        ������������������������       �                     @        K       L                 0c@z�G�z�?             @        ������������������������       �                     @        M       N                 p�w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        Q       R                 03k:@x��}�?            �K@        ������������������������       �                      @        S       n                   �J@ {��e�?            �J@       T       m                   �H@�%^�?            �E@       U       ^                   �<@:�&���?            �C@        V       ]                     �?�z�G��?             $@       W       X                 `ffC@և���X�?             @        ������������������������       �                      @        Y       Z                    7@z�G�z�?             @        ������������������������       �                      @        [       \                 ��I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        _       `                 �|Y>@\-��p�?             =@        ������������������������       �                     ,@        a       h                   �E@������?	             .@        b       g                   �C@      �?             @       c       f                    A@      �?             @       d       e                   @K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        i       j                    �?�����H�?             "@        ������������������������       �                     �?        k       l                 03C@@      �?              @        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        p       w                 @�:x@     ��?             @@       q       r                 0w�W@`Jj��?             ?@       ������������������������       �                     4@        s       t                    �?"pc�
�?             &@        ������������������������       �                     @        u       v                    6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        y       �                    �?������?�            w@        z       �                    �?Z�K�D��?;            �W@        {       |                 ���@П[;U��?             =@        ������������������������       �                     @        }       �                 �&�)@��H�}�?             9@       ~                           �?@4և���?             ,@        ������������������������       �                      @        �       �                    �?�8��8��?
             (@       ������������������������       �        	             &@        ������������������������       �                     �?        �       �                 �?�-@���!pc�?             &@       �       �                   �0@      �?              @        �       �                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @C@
��[��?(            @P@       �       �                   �>@��N`.�?#            �K@       �       �                   �0@ �o_��?             I@        ������������������������       �                     @        �       �                 P�@f.i��n�?            �F@        �       �                 pf�@      �?              @        ������������������������       �                     @        �       �                 �&B@      �?             @       �       �                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 03�0@��G���?            �B@       �       �                    �?�q�q�?             8@       �       �                    �?��s����?             5@       �       �                 �|�;@r�q��?	             2@       ������������������������       �                     (@        �       �                 pf&(@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �&@�q�q�?             @        ������������������������       �                     �?        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        �       �                   @B@z�G�z�?             @        ������������������������       �                     @        �       �                 ��|4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?䦳	�R�?�            0q@       �       �                 ��q1@`U���H�?�            �n@       �       �                    ,@���^���?�            �l@        ������������������������       �                     �?        �       �                    �?��8"W�?�            �l@        �       �                   �6@     ��?             @@        �       �                 ��y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|Y=@XB���?             =@        �       �                   @@      �?             @        ������������������������       �                      @        �       �                 ��Y&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     9@        �       �                   @@@TE½I�?{            �h@       �       �                    �?l{��b��?e            �c@        �       �                 �|Y=@$�q-�?             :@        �       �                  ��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���@�nkK�?             7@        ������������������������       �                      @        �       �                   @'@��S�ۿ?	             .@       ������������������������       �$�q-�?             *@        ������������������������       �                      @        �       �                 �?�@�U�=���?V            �`@        �       �                   �7@���N8�?*            �O@        ������������������������       �                     <@        �       �                   �8@�#-���?            �A@        �       �                 `fF@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�<@ 	��p�?             =@        ������������������������       �        	             &@        �       �                  sW@�����H�?             2@        �       �                 pf�@      �?              @        ������������������������       �                     @        �       �                 �|Y>@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 0SE @�θV�?,            @Q@        �       �                    3@r�q��?             >@        ������������������������       �                      @        �       �                    ?@ �Cc}�?             <@       �       �                   �4@�>����?             ;@        �       �                 @3�@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                 �|Y=@���7�?             6@        ������������������������       �                     @        �       �                 �|�=@      �?
             0@       �       �                 ��) @@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|�=@�7��?            �C@       ������������������������       �                    �A@        �       �                 ��Y)@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �C@        �       �                    ;@�q�q�?             .@        ������������������������       �                     @        �       �                 �|�<@      �?              @        ������������������������       �                      @        �       �                 �T)D@      �?             @       �       �                 X�,A@      �?             @       �       �                 м�5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?z�G�z�?             >@        �       �                   �2@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������T1�m��?X�]$���?*�Y7�"�?v�)�Y7�?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        vշ����?U��
R�?�>��x�?�ƃ�D�?�~j�t��?X9��v�?�E(B�?��^����?ہ�v`��?�3J���?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?        ^Cy�5�?(������?�$I�$I�?۶m۶m�?�$I�$I�?�m۶m��?              �?      �?                      �?�������?�������?              �?      �?      �?      �?                      �?              �?�-؂-��?�I��I��?��g�`�?�g�`�|�?�������?�?      �?        ��}��}�?AA�?      �?              �?      �?      �?        GX�i���?�{a���?�?�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?              �?      �?�p=
ף�?���Q��?�������?333333�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?              �?      �?      �?      �?              �?      �?              �?      �?        �������?�������?              �?�������?�������?              �?      �?      �?      �?                      �?      �?        pX���o�?A��)A�?              �?~�	�[�?
�[���?�}A_��?�}A_�?�A�A�?�o��o��?ffffff�?333333�?�$I�$I�?۶m۶m�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        a����?�{a���?      �?        wwwwww�?�?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�q�q�?�q�q�?      �?              �?      �?�������?�������?      �?                      �?      �?              �?      �?���{��?�B!��?      �?        /�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?G:l��F�?�On���?R�٨�l�?]AL� &�?��=���?�{a���?      �?        
ףp=
�?{�G�z�?�$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?t�E]t�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?7r#7r#�?�����?��oX���?� O	��?
ףp=
�?�Q����?      �?        �`�`�?�>�>��?      �?      �?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?#�u�)��?v�)�Y7�?�������?�������?z��y���?�a�a�?�������?UUUUUU�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        �������?�������?              �?      �?      �?      �?                      �?      �?        G�kĿF�?���ʽ?�[���?d �?�*�?ܯK*��?���ϱ?              �?b��g��?�G�İ?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?GX�i���?�{a���?      �?      �?      �?              �?      �?              �?      �?              �?        �wT���?&���0�?${�ґ�?�&��jq�?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?                      �?�Mozӛ�?d!Y�B�?      �?        �������?�?�؉�؉�?;�;��?      �?        �M6�d��?e�M6�d�?��y��y�?�a�a�?      �?        �A�A�?_�_�?�������?UUUUUU�?              �?      �?        ������?�{a���?      �?        �q�q�?�q�q�?      �?      �?      �?        333333�?�������?      �?      �?      �?              �?        ̵s���?�Q�g���?�������?UUUUUU�?              �?%I�$I��?۶m۶m�?�Kh/��?h/�����?�������?�������?      �?      �?      �?        �.�袋�?F]t�E�?      �?              �?      �?n۶m۶�?�$I�$I�?      �?                      �?      �?                      �?��[��[�?�A�A�?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?      �?      �?      �?      �?                      �?      �?                      �?�������?�������?�$I�$I�?۶m۶m�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ\bshG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                  x#J@���%&�?�           8�@              [                 `f�%@^djJ��?k           �@                                   �?C؇eY�?�            �p@                                  �0@�q�q�?-            @Q@        ������������������������       �                     @                                   �?     ��?)             P@                                ���@�����?
             3@        ������������������������       �                     @        	       
                    �?     ��?	             0@       ������������������������       �                     *@        ������������������������       �                     @                                �|Y=@�����H�?            �F@                                   �?�q�q�?             (@                                  ;@���Q��?             $@                               ���@      �?              @        ������������������������       �                     @                                  �2@      �?             @        ������������������������       �                     �?                                  �5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                   ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �@@               0                    �?`{��T��?            @i@                                  �3@���Q��?            �A@                                �&B@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                %                 P�@�q�q�?             >@        !       $                 pff@؇���X�?             @        "       #                 �|�9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        &       +                 `f�$@�㙢�c�?             7@       '       *                 `��!@@4և���?             ,@       (       )                 `�X!@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ,       /                     @�q�q�?             "@       -       .                   �J@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        1       >                   �<@ eD5�Ҽ?j            �d@        2       =                   �3@��pBI�?/            @R@        3       4                   �1@���}<S�?             7@        ������������������������       �                     @        5       :                   �2@�t����?
             1@        6       7                 ��@؇���X�?             @        ������������������������       �                     @        8       9                 ��Y @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ;       <                     @ףp=
�?             $@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �        !             I@        ?       N                 ��) @dP-���?;            �W@       @       A                 ��@�7��?0            �S@        ������������������������       �                     >@        B       E                 �|�>@�8��8��?             H@       C       D                 ��L@Pa�	�?            �@@        ������������������������       ��q�q�?             @        ������������������������       �                     >@        F       M                 @3�@z�G�z�?             .@       G       L                   �C@�q�q�?             "@       H       I                 �?�@      �?             @        ������������������������       �                      @        J       K                   �A@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        O       P                 ��y @      �?             0@        ������������������������       �                      @        Q       R                     @؇���X�?
             ,@        ������������������������       �                     @        S       Z                    ?@z�G�z�?             $@        T       U                 ���"@      �?             @        ������������������������       �                     �?        V       W                 �|Y=@�q�q�?             @        ������������������������       �                     �?        X       Y                 �|�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        \       �                     @��c�o��?�            0s@       ]       �                    �?�-�c��?r            �f@       ^       �                 0��I@*O���?X             b@       _       �                  �>I@F�����?S            �`@       `                        03�9@p�ݯ��?R            �`@        a       n                    �?����S��?%             M@        b       c                    �?�t����?             1@        ������������������������       �                     @        d       m                   �*@r�q��?	             (@       e       f                 `f�)@      �?              @        ������������������������       �                     �?        g       h                    :@����X�?             @        ������������������������       �                     �?        i       j                   �A@r�q��?             @       ������������������������       �                     @        k       l                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        o       p                     �?������?            �D@        ������������������������       �                      @        q       r                 �|Y=@�7��?            �C@        ������������������������       �        
             2@        s       v                 �|Y?@�����?             5@        t       u                 ��,@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        w       ~                   @F@�X�<ݺ?             2@       x       y                   �)@      �?              @        ������������������������       �                      @        z       }                    1@r�q��?             @       {       |                   @D@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?v�(��O�?-            �R@        �       �                    �?�X�<ݺ?             2@        �       �                 ��A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             ,@        �       �                 ��$:@�d�����?!            �L@        ������������������������       �        	             2@        �       �                  �>@�n_Y�K�?            �C@       �       �                    �?� �	��?             9@        �       �                 �ܵ<@z�G�z�?             @        �       �                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �=@      �?             4@       �       �                    J@      �?	             0@       �       �                    D@      �?              @        ������������������������       �                     @        �       �                   `G@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    C@@4և���?	             ,@       ������������������������       �                     $@        �       �                    H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�?�'�@�?             C@        �       �                     �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �A@�FVQ&�?            �@@       �       �                   �(@(;L]n�?             >@        ������������������������       �                     �?        ������������������������       �                     =@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?J��	�y�?M            @_@        �       �                 03�7@�G\�c�?&            @P@       �       �                   �:@؀�:M�?            �B@        �       �                    �?      �?             0@        �       �                    �?և���X�?             @       �       �                   �-@���Q��?             @       �       �                 �&�)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�<ݚ�?             "@       �       �                   @1@      �?              @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��.@��s����?             5@        �       �                    �?X�<ݚ�?             "@       �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?؇���X�?             <@        ������������������������       �                     �?        �       �                    @�����H�?             ;@        �       �                    �?؇���X�?             ,@        ������������������������       �                      @        �       �                    @r�q��?             (@        �       �                    @�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @$�q-�?             *@        ������������������������       �                      @        �       �                   @C@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 ��*@z�G�z�?'             N@        ������������������������       �                     @        �       �                 �J/@؇���X�?$             L@        ������������������������       �        	             0@        �       �                    �?z�G�z�?             D@        �       �                 03�6@�S����?             3@       ������������������������       �                     (@        �       �                 03�7@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @���N8�?             5@        ������������������������       �                     @        �       �                    0@     ��?             0@        ������������������������       �                     @        �       �                    @�8��8��?
             (@        ������������������������       �                     �?        ������������������������       �        	             &@        �       �                    �?x%[VY[�?Q            �`@       �       �                 ���Q@ĴF���?2            �T@        �       �                 �|�=@r�q��?             >@       �       �                     @     ��?	             0@       ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     ,@        �       �                    "@ ��WV�?"             J@        ������������������������       �                      @        ������������������������       �        !             I@        �       �                    �?��.k���?            �I@        �       �                 ��UO@���Q��?             4@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                 p"�X@����X�?	             ,@        ������������������������       �                     @        �       �                 @�ys@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �                          �;@���@M^�?             ?@        �       �                 0wkS@z�G�z�?             $@       �       �                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                              �|Y>@��s����?             5@        ������������������������       �                     @                                 A@������?
             .@        ������������������������       �                      @                              03�U@8�Z$���?	             *@       ������������������������       �                      @              
                  �L@���Q��?             @             	                ���a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������g *��?�0���M�?�.Lj��?�g+��?%��J?s�?m�}�3�?UUUUUU�?UUUUUU�?              �?      �?      �?^Cy�5�?Q^Cy��?      �?              �?      �?              �?      �?        �q�q�?�q�q�?�������?�������?333333�?�������?      �?      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?      �?        !w�l�2�?�F�tj�?333333�?�������?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?�7��Mo�?d!Y�B�?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?      �?                      �?      �?        UUUUUU�?UUUUUU�?�������?333333�?              �?      �?              �?        :�2	v�?\��l���?���Ǐ�?����?ӛ���7�?d!Y�B�?      �?        <<<<<<�?�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?        �����F�?W�+�ɵ?��[��[�?�A�A�?      �?        UUUUUU�?UUUUUU�?|���?|���?UUUUUU�?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        �)��-�?��F���?���?>��=���?�q�q�?�q�q�?�>�>��?؂-؂-�?^Cy�5�?Cy�5��?X�i���?O#,�4��?�?<<<<<<�?              �?UUUUUU�?�������?      �?      �?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?p>�cp�?������?      �?        ��[��[�?�A�A�?      �?        =��<���?�a�a�?UUUUUU�?UUUUUU�?              �?      �?        ��8��8�?�q�q�?      �?      �?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?              �?        Y�%�X�?O贁N�?�q�q�?��8��8�?      �?      �?      �?                      �?              �?Cy�5��?y�5���?      �?        ;�;��?ى�؉��?)\���(�?�Q����?�������?�������?      �?      �?      �?                      �?              �?      �?      �?      �?      �?      �?      �?              �?      �?      �?      �?                      �?      �?                      �?n۶m۶�?�$I�$I�?      �?              �?      �?              �?      �?                      �?�q�q�?�q�q�?              �?      �?        y�5���?������?333333�?�������?      �?                      �?|���?>����?�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        j�t��?+�����?S+�R+��?[��Z���?v�)�Y7�?E>�S��?      �?      �?۶m۶m�?�$I�$I�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?        9��8���?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�a�a�?z��y���?�q�q�?r�q��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?۶m۶m�?�$I�$I�?              �?�q�q�?�q�q�?۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �؉�؉�?;�;��?      �?        ]t�E�?F]t�E�?              �?      �?        �������?�������?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?(������?^Cy�5�?      �?        �$I�$I�?۶m۶m�?              �?      �?        �a�a�?��y��y�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �d\�?}s����?ە�]�ڵ?E�JԮD�?UUUUUU�?�������?      �?      �?              �?      �?                      �?;�;��?O��N���?      �?                      �?�������?�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?�m۶m��?              �?�$I�$I�?۶m۶m�?      �?                      �?�s�9��?�c�1��?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?z��y���?�a�a�?      �?        wwwwww�?�?              �?;�;��?;�;��?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0Kh2h3h4hph<�h=Kub��������                           @ʡ�;S��?�           8�@                                    @�4F����?            �D@        ������������������������       �        	             (@                                ��|2@П[;U��?             =@        ������������������������       �                     &@                                   @�E��ӭ�?             2@        ������������������������       �                     "@               	                    �?X�<ݚ�?             "@        ������������������������       �                      @        
                           �?����X�?             @                               `f�:@z�G�z�?             @        ������������������������       �                     @                                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               Z                    �?�b�]�?�           ��@               +                     @(����?�            `l@              $                   �B@���}��?L            �`@              #                   �;@��:x�ٳ?7            �X@                                    �?���}<S�?             G@        ������������������������       �                     6@                                   �9@r�q��?             8@                                 �+@P���Q�?             4@                                   �?      �?             @        ������������������������       �                     �?                                  �6@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        !       "                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �J@        %       &                   @C@�t����?             A@        ������������������������       �                      @        '       *                    �?      �?             @@        (       )                 83F@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     3@        ,       Y                   �@@��V�I��?=            �W@       -       L                    �?�p ��?5            �T@       .       ;                    �?�q�q�?#             H@       /       6                    �?�r����?             >@        0       1                 H�%@�z�G��?             $@        ������������������������       �                     @        2       5                 ���,@���Q��?             @       3       4                   �-@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        7       8                 �|�9@P���Q�?             4@        ������������������������       �                     @        9       :                  ��@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �        
             *@        <       E                   �9@�q�q�?             2@       =       >                 pf�@�θ�?
             *@        ������������������������       �                      @        ?       D                    3@�C��2(�?             &@        @       A                 ��!@z�G�z�?             @        ������������������������       �                      @        B       C                 `F�+@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        F       G                 @3�@���Q��?             @        ������������������������       �                     �?        H       I                 @3�,@      �?             @        ������������������������       �                      @        J       K                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        M       X                 ��l4@�t����?             A@       N       W                 �|Y=@      �?
             4@       O       P                   �#@�q�q�?             .@        ������������������������       �                     @        Q       R                    5@�eP*L��?             &@        ������������������������       �                     @        S       T                    <@؇���X�?             @        ������������������������       �                     @        U       V                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     (@        [       �                     �?��:�Xn�?           �{@        \       �                    �?�q�q�?=             X@       ]       d                   �<@�H�a��?5            @U@        ^       _                 `f�D@�	j*D�?             *@        ������������������������       �                     @        `       a                    6@      �?              @        ������������������������       �                      @        b       c                   �:@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        e       n                    �?      �?-             R@        f       g                   @@@      �?             4@        ������������������������       �                     @        h       m                   �H@�n_Y�K�?	             *@       i       l                  xCH@r�q��?             @        j       k                   �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        o       �                   @J@      �?              J@       p       �                   �G@�����?             C@       q       �                   �F@�'�`d�?            �@@       r       y                   �>@      �?             <@        s       t                 �|Y=@�q�q�?	             (@        ������������������������       �                      @        u       v                 �̌/@      �?             $@        ������������������������       �                     @        w       x                   �C@r�q��?             @       ������������������������       �                     @        ������������������������       �      �?              @        z       {                 `f�K@      �?	             0@       ������������������������       �                     &@        |       }                 �|Y>@���Q��?             @        ������������������������       �                      @        ~                        03�Q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 `fF<@@4և���?             ,@        ������������������������       �                      @        �       �                  )?@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �4@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    @@���މ�?�            �u@       �       �                     @؇���X�?�            �p@        �       �                    &@Pa�	�?            �@@        �       �                    @ףp=
�?	             $@        ������������������������       �                     @        �       �                   �5@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        �       �                 �T�I@�Nx�1�?�             m@       �       �                    �?*
;&���?�            �l@        �       �                   �6@">�֕�?            �A@        �       �                   �2@      �?              @       �       �                 �x"@�q�q�?             @        ������������������������       �                     �?        �       �                 �y.@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|=@�+$�jP�?             ;@        ������������������������       �                     @        �       �                 �|�=@      �?             4@       �       �                    �?�E��ӭ�?             2@       �       �                 ���@�r����?
             .@        ������������������������       �                     @        �       �                   @@z�G�z�?             $@       ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                  ��@�?�<��?s            `h@        �       �                 ���@XB���?             =@        �       �                 ���@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �        
             1@        �       �                    �?�/ C-��?a            �d@       �       �                 �|�=@؇���X�?Z            @c@       �       �                   �<@L������?T            @b@       �       �                 0S5 @�7��?/            �S@       �       �                   �4@�:�^���?             �F@        �       �                   �3@�	j*D�?             *@       �       �                 pf�@      �?              @        ������������������������       �                      @        �       �                   �1@      �?             @        ������������������������       �      �?             @        ������������������������       �      �?              @        �       �                 P�@z�G�z�?             @        ������������������������       �                      @        �       �                 @3�@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @@        ������������������������       �                    �@@        �       �                 �|Y=@@�0�!��?%             Q@        �       �                   @@�q�q�?             "@        ������������������������       �                     @        �       �                 ���"@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 м�5@�j��b�?!            �M@       �       �                 �Y5@x�}b~|�?            �L@        �       �                 ��@d}h���?
             ,@       ������������������������       ��8��8��?	             (@        ������������������������       �                      @        �       �                    �? �#�Ѵ�?            �E@        ������������������������       �                     "@        �       �                 ��) @�IєX�?             A@       ������������������������       �                     7@        �       �                 �̜!@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �>@      �?              @        ������������������������       �                      @        �       �                   �?@�q�q�?             @        �       �                 pff@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 P�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        �       �                 �̌4@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @ �)���?5            @T@        �       �                   @A@      �?             @@        �       �                    1@؇���X�?             @        �       �                 `fF)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     9@        ������������������������       �                    �H@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������N���I5�?d�~`l��?KԮD�J�?ە�]���?              �?��=���?�{a���?              �?�q�q�?r�q��?      �?        �q�q�?r�q��?      �?        �$I�$I�?�m۶m��?�������?�������?              �?      �?      �?              �?      �?              �?      �?              �?      �?        �������?�R,Z�?�D�����?�]/����?���̮?4�τ?�?[�R�֯�?
�����?d!Y�B�?ӛ���7�?              �?UUUUUU�?�������?�������?ffffff�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?                      �?�?<<<<<<�?      �?              �?      �?;�;��?;�;��?      �?                      �?              �?G}g����?r1����?8��18�?dp>�c�?UUUUUU�?UUUUUU�?�?�������?333333�?ffffff�?              �?333333�?�������?      �?      �?      �?                      �?      �?        �������?ffffff�?              �?�$I�$I�?n۶m۶�?      �?                      �?UUUUUU�?UUUUUU�?ى�؉��?�؉�؉�?              �?]t�E�?F]t�E�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �������?333333�?      �?              �?      �?              �?      �?      �?      �?                      �?�������?�������?      �?      �?UUUUUU�?UUUUUU�?              �?]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?              �?              �?              �?        �-�)�?�cI��[�?�������?�������?�������?TTTTTT�?;�;��?vb'vb'�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?      �?        ;�;��?ى�؉��?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?              �?      �?Q^Cy��?^Cy�5�?6�d�M6�?'�l��&�?      �?      �?�������?�������?      �?              �?      �?      �?        UUUUUU�?�������?              �?      �?      �?      �?      �?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?n۶m۶�?�$I�$I�?      �?        �������?UUUUUU�?              �?      �?        ]t�E�?F]t�E�?              �?      �?        <=�	Ig�?"F��ż?۶m۶m�?�$I�$I�?|���?|���?�������?�������?      �?        �������?�������?              �?      �?              �?        �X����?����S�?���,d!�?8��Moz�?_�_��?�A�A�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?/�����?B{	�%��?      �?              �?      �?�q�q�?r�q��?�������?�?      �?        �������?�������?�m۶m��?�$I�$I�?      �?                      �?      �?        �����? �����?GX�i���?�{a���?UUUUUU�?UUUUUU�?      �?                      �?      �?        8�:����?"�%��?۶m۶m�?�$I�$I�?�Ǐ?~�?����?��[��[�?�A�A�?}�'}�'�?l�l��?vb'vb'�?;�;��?      �?      �?      �?              �?      �?      �?      �?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?              �?        ZZZZZZ�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�N��?��/���?�YLg1�?Lg1��t�?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?              �?�/����?�}A_Ч?      �?        �?�?      �?        /�袋.�?F]t�E�?              �?      �?              �?      �?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?X�<ݚ�?�����H�?      �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJj�c;hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������       b                     @|��;;��?�           8�@               S                    �?ޣ]M��?�            �t@              ,                     �?n�QJ���?�            `o@                                  �?և���X�?X            �a@        ������������������������       �        %            �K@               %                   @J@�t����?3            @U@                               03:@:PZ(8?�?,            @R@        ������������������������       �                     @        	       $                   �G@�T��5m�?(            �P@       
       #                   �E@V��z4�?%             O@                                 @@@��C���?            �G@                                  �?������?             A@                                `ffA@؇���X�?             ,@                                ���<@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                  �<@�z�G��?             4@                                `f&F@�q�q�?             @       ������������������������       �                     @                                   7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  �>@؇���X�?
             ,@                                �|Y=@      �?             @        ������������������������       �                     �?                                `fF<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@                                 `�iJ@8�Z$���?             *@       ������������������������       �                     @        !       "                 03�Q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     @        &       '                    �?�8��8��?             (@        ������������������������       �                     @        (       )                 `fF<@      �?              @        ������������������������       �                     @        *       +                   �?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        -       >                    �?���I���?E            �[@        .       =                 ��*@�8��8��?             B@       /       <                   �J@ȵHPS!�?             :@       0       5                   �9@HP�s��?             9@        1       2                    �?z�G�z�?             @        ������������������������       �                      @        3       4                   �6@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        6       7                    �?P���Q�?             4@        ������������������������       �                      @        8       9                   �'@�X�<ݺ?             2@        ������������������������       �                     "@        :       ;                   �B@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ?       @                    �?��S�ۿ?-            �R@        ������������������������       �                     @        A       H                   �@@����p�?(             Q@       B       G                    &@������?             B@        C       D                    @�C��2(�?	             &@        ������������������������       �                     @        E       F                    5@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     9@        I       J                   @A@      �?             @@        ������������������������       �                     @        K       L                 `f�)@XB���?             =@        ������������������������       �                     "@        M       R                   �*@P���Q�?             4@       N       Q                   �F@�8��8��?             (@        O       P                   @D@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        T       W                    �?��مD�?3            @S@       U       V                    @`'�J�?            �I@        ������������������������       �                      @        ������������������������       �                    �H@        X       ]                   �7@
j*D>�?             :@        Y       Z                    4@ףp=
�?	             $@       ������������������������       �                     @        [       \                 `�B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ^       a                    �?      �?             0@       _       `                 �̾w@؇���X�?	             ,@       ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                      @        c       p                    @��<f*�?�            �w@        d       e                    �?���N8�?             5@        ������������������������       �                     @        f       g                    �?�E��ӭ�?             2@        ������������������������       �                     @        h       k                    �?�eP*L��?             &@        i       j                    @      �?             @        ������������������������       �                     @        ������������������������       �                     @        l       o                    @���Q��?             @       m       n                 pf�C@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        q       �                    �?~_d+�^�?�            �v@        r       �                   @B@��7 ���??            �W@       s       �                 `v�6@�!>�R�?9            �T@       t       {                 �̌@|�U&k�?3            �R@        u       z                 ���@�nkK�?             7@        v       w                 �|Y:@z�G�z�?             @       ������������������������       �                     @        x       y                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        |       �                 pF�%@�~8�e�?"            �I@        }       �                    �?�	j*D�?
             *@       ~                           �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �7@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �*@P����?             C@        ������������������������       �                     "@        �       �                 �?�-@П[;U��?             =@        �       �                 ���,@؇���X�?             @       �       �                   �-@z�G�z�?             @        ������������������������       �                      @        �       �                   �0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�X����?             6@        �       �                 �|Y=@؇���X�?             @        ������������������������       �                      @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���Q��?
             .@       �       �                 ���1@��
ц��?	             *@       �       �                 �|�;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                     @        �       �                 ���4@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     &@        �       �                   @@@��v����?�            �p@       �       �                    �?�MI8d�?�            �k@        �       �                 ���@     ��?             @@        �       �                 ��y@�C��2(�?             &@        ������������������������       �                     @        �       �                 �|�9@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    7@�ՙ/�?             5@        �       �                   �2@���Q��?             $@       �       �                    -@�q�q�?             @       �       �                    '@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?"pc�
�?             &@       �       �                 �|Y=@ףp=
�?             $@        �       �                   �;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��,�5�?s            �g@        �       �                 ���@�חF�P�?             ?@        ������������������������       �                     @        �       �                 ��(@z�G�z�?             9@       �       �                 �|Y=@�	j*D�?             *@        ������������������������       �                      @        ������������������������       �"pc�
�?             &@        �       �                 �|�2@�8��8��?             (@        ������������������������       �                     @        �       �                   `3@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�S�%3��?`            �c@       �       �                   �>@̻L&��?Z            �b@       �       �                   �7@��ׄ��?T            `a@        �       �                   �0@ ������?$            �O@        �       �                 pFD!@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      M@        �       �                 ��) @�S����?0             S@       �       �                   @8@      �?"             H@        �       �                 `fF@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��L@���7�?             F@        �       �                 �|Y=@"pc�
�?             &@        ������������������������       �                     @        �       �                 ��,@      �?              @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                    �@@        �       �                   �<@��X��?             <@       �       �                   �;@     ��?             0@        �       �                   �:@և���X�?             @       �       �                 �T)D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                 �|�=@      �?             (@       �       �                 `��!@�eP*L��?             &@        ������������������������       �                      @        �       �                 �|Y=@�q�q�?             "@        �       �                 ���"@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �&B@      �?             (@        ������������������������       �                     �?        �       �                   �?@"pc�
�?             &@        ������������������������       �                     @        �       �                 P�@      �?              @        ������������������������       �                      @        �       �                 d�@@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     G@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������|d�_Z�?�7s@K�?E�JԮD�?^�ڕ�]�?������?���0p�?۶m۶m�?�$I�$I�?              �?�������?�������?�W�^�z�?�P�B�
�?      �?        9��_���?���@���?2�c�1�?�s�9��?L� &W�?g���Q��?xxxxxx�?�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ffffff�?333333�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?      �?              �?      �?        �Ps��?�^����?UUUUUU�?UUUUUU�?�؉�؉�?��N��N�?{�G�z�?q=
ףp�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?ffffff�?              �?�q�q�?��8��8�?              �?�q�q�?�q�q�?              �?      �?              �?                      �?�������?�?      �?        �������?�����Ҳ?�q�q�?�q�q�?]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?              �?      �?              �?GX�i���?�{a���?      �?        ffffff�?�������?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?      �?              �?        �	qV~B�?��cj`��?�?�������?      �?                      �?b'vb'v�?;�;��?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?۶m۶m�?�$I�$I�?      �?                      �?      �?        �����d�?�
$6�?��y��y�?�a�a�?              �?r�q��?�q�q�?              �?]t�E�?t�E]t�?      �?      �?      �?                      �?�������?333333�?      �?      �?              �?      �?              �?        ��T4O�?�o��.��?�����F�?1���\�?��k���?+Jx���?E>�S��?�`�|��?d!Y�B�?�Mozӛ�?�������?�������?              �?      �?      �?              �?      �?                      �?�������?222222�?vb'vb'�?;�;��?�q�q�?�q�q�?              �?      �?              �?      �?              �?      �?        Q^Cy��?�P^Cy�?              �?��=���?�{a���?۶m۶m�?�$I�$I�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ]t�E]�?�E]t��?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?        �������?333333�?�؉�؉�?�;�;�?UUUUUU�?�������?      �?                      �?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?                      �?      �?              �?        5&����?*g��1�?��L���?L�Ϻ��?      �?      �?]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        �<��<��?�a�a�?�������?333333�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?/�袋.�?F]t�E�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?>�ĩ�s�?#�X�0�?�Zk����?��RJ)��?      �?        �������?�������?vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?      �?                      �?T�p���?�.=���?�Y�vV�?��JL%��?�Ke{��?��$D�?��}��}�?AA�?�������?�������?      �?      �?      �?              �?        (������?^Cy�5�?      �?      �?      �?      �?              �?      �?        �.�袋�?F]t�E�?/�袋.�?F]t�E�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?        n۶m۶�?%I�$I��?      �?      �?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?      �?              �?      �?t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?      �?      �?      �?        F]t�E�?/�袋.�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJGԙGhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM+hjh))��}�(h,h/h0M+��h2h3h4hph<�h=Kub������       b                    �?e�L��?�           8�@                                   (@n���C�?�             n@               
                    @��
ц��?             :@                               03�=@������?             .@       ������������������������       �                     "@                                     @�q�q�?             @        ������������������������       �                      @               	                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @                                03;@�C��2(�?             &@                                   @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               %                     @7���?�            �j@                                   �?P#aE�?M            �`@                                 �H@��v$���?(            �N@       ������������������������       �                      J@                                �DD@�����H�?             "@                                ���;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               $                    �?�n���?%             R@                               ���&@�q��/��?             G@                                  �J@�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @               #                   �;@�FVQ&�?            �@@                                    �?�q�q�?             @        ������������������������       �                      @        !       "                   �5@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ;@        ������������������������       �                     :@        &       [                   �A@�Je\���?7            @T@       '       D                 �|Y=@Pa�.l�?0            �P@       (       7                   �6@      �?             B@       )       2                 ��,#@p�ݯ��?             3@       *       1                   �3@8�Z$���?             *@        +       ,                    �?����X�?             @        ������������������������       �                     �?        -       .                   �1@�q�q�?             @        ������������������������       �                      @        /       0                   !@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        3       6                    3@r�q��?             @       4       5                 �K(@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        8       =                   �&@ҳ�wY;�?             1@       9       <                 P�@ףp=
�?             $@        :       ;                   �9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        >       C                   �;@����X�?             @       ?       @                    9@r�q��?             @        ������������������������       �                     @        A       B                 @3�,@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        E       Z                 ��Y7@f���M�?             ?@       F       K                  ��@�θ�?             :@        G       H                    �?$�q-�?	             *@        ������������������������       �                      @        I       J                 ���@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        L       Y                    @@�n_Y�K�?
             *@       M       X                 03C3@�q�q�?	             (@       N       W                    �?����X�?             @       O       V                   �0@�q�q�?             @       P       Q                 ��� @      �?             @        ������������������������       �                     �?        R       S                 �?$'@�q�q�?             @        ������������������������       �                     �?        T       U                  S�-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        \       ]                 ��A>@؇���X�?             ,@       ������������������������       �                     $@        ^       a                    @      �?             @       _       `                   �C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        c       �                     �?�p�ҝ�?,           p}@        d       e                 ��$:@*Mp����?E            �Y@        ������������������������       �                     &@        f       �                    �?�n_Y�K�?>            �V@       g       ~                  �>@�!�,�E�?3            @R@        h       }                    K@����"�?             =@       i       n                    �?��<b���?             7@        j       k                 �|�=@z�G�z�?             @        ������������������������       �                      @        l       m                   @@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        o       p                 03k:@�<ݚ�?             2@        ������������������������       �                     @        q       r                 �|Y=@������?
             .@        ������������������������       �                     �?        s       |                   `G@d}h���?	             ,@       t       {                   �F@���!pc�?             &@       u       x                 �|�?@z�G�z�?             $@        v       w                 `fF<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        y       z                   �C@r�q��?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               �                  x#J@v�X��?             F@        �       �                 �|�<@�KM�]�?             3@        ������������������������       �                     �?        �       �                    �?�X�<ݺ?             2@        �       �                 `f�A@      �?              @        �       �                 X�lA@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �8@� �	��?             9@        ������������������������       �                     @        �       �                    <@�G�z��?             4@        ������������������������       �                     @        �       �                    �?�	j*D�?             *@        �       �                 �UkT@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �B@���!pc�?	             &@        ������������������������       �                     @        �       �                   �E@      �?              @        ������������������������       �                      @        �       �                    H@r�q��?             @        ������������������������       �                     @        �       �                 ���W@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�<ݚ�?             2@       �       �                   @B@������?             .@        �       �                   �?@�q�q�?             @       �       �                 ��-a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �       �                    �?�p ��?�            w@        �       �                 ��i @R�}e�.�?             J@       �       �                    �?��a�n`�?             ?@       �       �                 ���@ףp=
�?             >@        �       �                 03S@؇���X�?             ,@        ������������������������       �                     �?        �       �                 �|�9@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        �       �                 �|Y=@      �?	             0@        �       �                   @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     �?        �       �                     @�G��l��?
             5@        �       �                 `��.@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    /@�	j*D�?             *@        �       �                 =
�@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 03�-@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @ ���:�?�            �s@        �       �                    �?$��$�L�?3            �S@       �       �                   �*@hA� �?,            �Q@       �       �                 `f�)@=QcG��?             �G@       �       �                    4@h�����?             <@        �       �                   �2@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     5@        �       �                   �A@�KM�]�?             3@       �       �                 �|Y;@      �?              @        ������������������������       �                     @        �       �                 �|�=@���Q��?             @        ������������������������       �                     �?        �       �                    @@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     &@        ������������������������       �                     7@        �       �                    :@X�<ݚ�?             "@        �       �                    *@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             @       �       �                   P@@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �?�@0y����?�            �m@        �       �                    �?0x�!���?D            �]@       �       �                    �?���U�?C            �\@        �       �                 �|Y=@@4և���?             <@        �       �                  ��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     9@        �       �                 �|Y=@ qP��B�?4            �U@       ������������������������       �                     I@        �       �                 pf�@�X�<ݺ?             B@        ������������������������       �                     1@        �       �                   �@�KM�]�?             3@        �       �                 �|Y>@�q�q�?             @        ������������������������       �                     �?        �       �                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     @        �                          �?������?T            �]@       �                         @@@V�a�� �?<            �U@       �                       м�5@�+e�X�?3            �R@       �       	                �|�=@"pc�
�?-            �P@       �       �                   �:@���5��?(            �L@        �       �                 pf� @$�q-�?             :@        �       �                   �4@z�G�z�?             $@       �       �                 @3�@���Q��?             @        ������������������������       �                     �?        �       �                   �1@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        �       �                    �?�חF�P�?             ?@        ������������������������       �                      @        �       �                   �;@д>��C�?             =@        ������������������������       �                     �?        �                        ��) @؇���X�?             <@        ������������������������       �                     &@                              pf� @������?
             1@        ������������������������       �                      @                              ���(@�r����?	             .@                              ���"@�q�q�?             @        ������������������������       �                     @                                �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        
                      ��Y)@X�<ݚ�?             "@                             ��l!@      �?              @                               �?@      �?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?                              03�7@�q�q�?             "@        ������������������������       �                      @                                 �?և���X�?             @        ������������������������       �                     �?                                 ;@�q�q�?             @        ������������������������       �                     @                              �|�>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             (@              *                   #@     ��?             @@             !                   @j���� �?             1@                                 �?z�G�z�?             @       ������������������������       �                     @                               pf�@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        "      %                   �?      �?             (@       #      $                   �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        &      '                `f�9@z�G�z�?             @        ������������������������       �                      @        (      )                ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        �*       h�h))��}�(h,h/h0M+KK��h2h3h4hVh<�h=Kub������������v�S(��?��X��?DDDDDD�?�������?�;�;�?�؉�؉�?�?wwwwww�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?]t�E�?F]t�E�?      �?      �?              �?      �?              �?        �@�Ե�?�/Ċ���?�qA��?�蛣o��?;ڼOqɐ?.�u�y�?              �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?r�qǱ?r�q��?��Mozӻ?�B����?�؉�؉�?ى�؉��?              �?      �?        |���?>����?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?              �?ԭ�a�2�?X�<ݚ�?5&����?��~5&�?      �?      �?Cy�5��?^Cy�5�?;�;��?;�;��?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?�������?UUUUUU�?      �?      �?              �?      �?              �?        �������?�������?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?�m۶m��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        ��Zk���?��RJ)��?�؉�؉�?ى�؉��?;�;��?�؉�؉�?              �?F]t�E�?]t�E�?      �?                      �?ى�؉��?;�;��?�������?�������?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?                      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �R��
��?�����/�?�?�������?      �?        ;�;��?ى�؉��?�&M�4i�?ٲe˖-�?�i��F�?	�=����?��Moz��?��,d!�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?9��8���?              �?�?wwwwww�?      �?        ۶m۶m�?I�$I�$�?t�E]t�?F]t�E�?�������?�������?      �?      �?      �?                      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        �.�袋�?颋.���?�k(���?(�����?              �?��8��8�?�q�q�?      �?      �?      �?      �?      �?                      �?      �?              �?        �Q����?)\���(�?      �?        �������?�������?              �?vb'vb'�?;�;��?      �?      �?              �?      �?        F]t�E�?t�E]t�?      �?              �?      �?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?9��8���?�q�q�?wwwwww�?�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        Q��+Q�?��+Q��?'vb'vb�?�;�;�?�s�9��?�c�1Ƹ?�������?�������?۶m۶m�?�$I�$I�?      �?        ;�;��?;�;��?              �?      �?              �?      �?      �?      �?      �?                      �?      �?              �?        ��y��y�?1�0��?      �?      �?              �?      �?        ;�;��?vb'vb'�?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?      �?                      �?�7W$O��?!�n�&�?��]-n��?�3���?���?_�_�?x6�;��?AL� &W�?�m۶m��?�$I�$I�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?        �k(���?(�����?      �?      �?      �?        333333�?�������?              �?      �?      �?      �?              �?      �?      �?              �?        �q�q�?r�q��?�������?�������?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�5�5�?��~���?�5�5�?	�#����?p�}��?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��}A�?�}A_З?      �?        ��8��8�?�q�q�?      �?        �k(���?(�����?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        xxxxxx�?�?��{a�?a���{�?R���Q�?���Q��?/�袋.�?F]t�E�?�}��?��Gp�?�؉�؉�?;�;��?�������?�������?333333�?�������?              �?      �?      �?      �?      �?      �?              �?              �?        �Zk����?��RJ)��?      �?        a���{�?|a���?              �?۶m۶m�?�$I�$I�?      �?        xxxxxx�?�?              �?�������?�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?r�q��?      �?      �?      �?      �?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?ZZZZZZ�?�������?�������?�������?      �?              �?      �?              �?      �?              �?      �?�$I�$I�?�m۶m��?      �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��AhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       b                 ���$@�4�O��?�           8�@                                ���@��j���?�            q@        ������������������������       �                     @@                                   �?�}�V���?�             n@                                   �?���@M^�?'             O@                                   �?     ��?             @@        ������������������������       �                     @               	                 ���@ܷ��?��?             =@        ������������������������       �                     &@        
                          �5@r�q��?             2@        ������������������������       �                      @                                  @@      �?
             0@                               �|=@      �?              @        ������������������������       �                      @                                �|�=@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                      @                                �|Y=@���Q��?             >@        ������������������������       �                     @                                   �?�q�����?             9@                               03@؇���X�?	             ,@                               ���@"pc�
�?             &@        ������������������������       �                     �?                                   �?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                 s�@�C��2(�?             &@        ������������������������       �                     @        ������������������������       �      �?              @                !                 ���@8�e����?o            `f@        ������������������������       �                      @        "       3                   �2@t���s��?n             f@        #       *                   �1@����X�?             5@       $       )                    �?d}h���?             ,@       %       (                 pf� @8�Z$���?             *@        &       '                 pf�@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        +       0                    �?և���X�?             @        ,       -                 P��@�q�q�?             @        ������������������������       �                     �?        .       /                 ��!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       2                 P��@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        4       a                   �C@�:�^���?`            �c@       5       `                   @C@�KM�]�?U            �`@       6       ?                    �?@v�禺�?T            �`@        7       8                   �3@��s����?             5@        ������������������������       �                     �?        9       >                 �|Y>@R���Q�?             4@       :       =                   �7@�KM�]�?
             3@        ;       <                 pff@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        @       S                 ��) @�L���?H            �[@       A       N                   �?@`��F:u�?7            �U@       B       I                 �?$@�g<a�?/            @S@        C       D                 ���@�IєX�?
             1@       ������������������������       �                     *@        E       H                 �|Y>@      �?             @       F       G                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        J       K                 @3�@ �.�?Ƞ?%             N@       ������������������������       �                     B@        L       M                   �3@ �q�q�?             8@        ������������������������       �      �?             @        ������������������������       �                     4@        O       R                   �@z�G�z�?             $@        P       Q                   @@@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        T       U                    9@�q�q�?             8@        ������������������������       �                     (@        V       _                   �?@�q�q�?	             (@       W       X                   �;@      �?              @        ������������������������       �                      @        Y       Z                   �<@      �?             @        ������������������������       �                      @        [       ^                 ��)"@      �?             @        \       ]                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     7@        c       �                     @#F���?           `{@       d       �                 `fFJ@�1:��?�            �r@       e       x                    �?.�����?u            @i@        f       w                    �?�:�^���?-            �S@       g       h                    �?      �?             L@        ������������������������       �                     @        i       j                     �?؇���X�?            �H@        ������������������������       �                     @        k       v                    L@���V��?            �F@       l       m                   �'@X�EQ]N�?            �E@        ������������������������       �                     "@        n       o                   �B@��hJ,�?             A@       ������������������������       �                     3@        p       q                   �C@�q�q�?             .@        ������������������������       �                     @        r       s                    5@r�q��?             (@       ������������������������       �                      @        t       u                   �E@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     6@        y       z                    #@��a�n`�?H             _@        ������������������������       �                     @        {       �                 ��D:@F�4�Dj�?E            �]@       |       �                   �*@������?+            �R@       }       ~                    �?r�q��?             H@        ������������������������       �                     @               �                 `f�)@:	��ʵ�?            �F@        �       �                    &@�C��2(�?             6@       �       �                    5@8�Z$���?             *@        ������������������������       ��q�q�?             @        ������������������������       �                     $@        ������������������������       �                     "@        �       �                    @@��+7��?             7@        ������������������������       �                     "@        �       �                   �A@և���X�?             ,@        ������������������������       �                     @        �       �                   @D@z�G�z�?             $@        ������������������������       �                     @        �       �                    G@�q�q�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     :@        �       �                   �R@�X����?             F@       �       �                     �?      �?             D@       �       �                  �>@:ɨ��?            �@@        �       �                    �?�θ�?	             *@        ������������������������       �                     @        �       �                   @=@�z�G��?             $@       �       �                   �F@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     4@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��.D��?A            @X@       �       �                 pf�Z@>a�����?!            �I@       �       �                    �? 	��p�?             =@       �       �                    �?$�q-�?             :@       ������������������������       �                     4@        �       �                    �?�q�q�?             @       ������������������������       �                     @        �       �                    F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?���!pc�?             6@       ������������������������       �        
             *@        �       �                 �̾w@�q�q�?             "@       �       �                   �1@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 03�M@���j��?              G@        ������������������������       �                      @        �       �                    �?P����?             C@       �       �                 ���a@�LQ�1	�?             7@       ������������������������       �        
             ,@        �       �                    �?�q�q�?             "@        ������������������������       �                     @        �       �                 Ъ�c@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                     �?�q�q�?
             .@       �       �                 �|�0@�n_Y�K�?             *@        ������������������������       �                     @        �       �                    J@�����H�?             "@       �       �                 ��#[@      �?             @        ������������������������       �                      @        �       �                  �6f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 pf�+@4V��X�?V            `a@        �       �                 `f�%@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �6@��O�;��?O             `@        �       �                 @3�4@"pc�
�?             �K@        �       �                    �?���|���?             6@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    '@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    $@p�ݯ��?	             3@        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?�FVQ&�?            �@@        ������������������������       �        	             1@        �       �                    �?      �?             0@       �       �                    @$�q-�?             *@        �       �                 ��T?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 ��T?@�q�q�?             @        ������������������������       �                     �?        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?4�B��?/            �R@        �       �                    �?��.k���?             A@        �       �                 X�l@@@4և���?             ,@       �       �                    �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �       �                    @R���Q�?             4@       �       �                    �?@�0�!��?             1@        �       �                  ��6@r�q��?             @        �       �                   �=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @34@"pc�
�?             &@        �       �                   �/@���Q��?             @       �       �                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �                          �?z�G�z�?             D@       �       	                   �?r֛w���?             ?@       �       �                   �:@R�}e�.�?             :@        �       �                 ��q1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �                       �|�>@R���Q�?             4@       �       �                 �|Y<@�t����?	             1@        ������������������������       �                     @        �       �                 м�5@؇���X�?             ,@       ������������������������       �                     "@                                  �?���Q��?             @                             03�7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                @B@�q�q�?             @                             �!B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        
                         �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������X�>�?2�N����?�������?Y�Y��?      �?        �a�a��?ynyn�?�s�9��?�c�1��?      �?      �?              �?��=���?a���{�?      �?        �������?UUUUUU�?              �?      �?      �?      �?      �?      �?        �������?UUUUUU�?      �?      �?      �?              �?        �������?333333�?              �?���Q��?�p=
ף�?�$I�$I�?۶m۶m�?F]t�E�?/�袋.�?              �?�������?�������?              �?      �?                      �?]t�E�?F]t�E�?      �?              �?      �?jr�y)�?�l|3�v�?              �?3��Yb�?k��2�?�m۶m��?�$I�$I�?I�$I�$�?۶m۶m�?;�;��?;�;��?333333�?�������?      �?                      �?      �?                      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?      �?                      �?� � �?�o��o��?�k(���?(�����?�d�M6��?6�d�M6�?z��y���?�a�a�?              �?333333�?333333�?�k(���?(�����?9��8���?�q�q�?              �?      �?              �?                      �?}���g�?L�Ϻ��?�u�7[��?Ȥx�L��?���8+�?�cj`?�?�?      �?              �?      �?      �?      �?      �?                      �?      �?        wwwwww�?�?      �?        �������?UUUUUU�?      �?      �?      �?        �������?�������?      �?      �?              �?      �?              �?        UUUUUU�?�������?      �?        �������?�������?      �?      �?              �?      �?      �?      �?              �?      �?      �?      �?              �?      �?                      �?      �?                      �?      �?        +���?�������?���̳��?������?h���Q�?0��<�]�?�o��o��?� � �?      �?      �?              �?�$I�$I�?۶m۶m�?              �?�>�>��?[�[��?qG�wĽ?w�qG�?              �?�������?KKKKKK�?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?              �?                      �?�c�1��?�s�9��?              �?��/���?�A�I��?��g�`��?к����?�������?UUUUUU�?      �?        ��O��O�?l�l��?]t�E�?F]t�E�?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?              �?        zӛ����?Y�B��?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        �E]t��?]t�E]�?      �?      �?N6�d�M�?e�M6�d�?�؉�؉�?ى�؉��?              �?333333�?ffffff�?۶m۶m�?�$I�$I�?              �?      �?                      �?      �?              �?                      �?��Id��?���fy�?�?�������?�{a���?������?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?t�E]t�?F]t�E�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?!Y�B�?ozӛ���?              �?Q^Cy��?�P^Cy�?Y�B��?��Moz��?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?;�;��?ى�؉��?              �?�q�q�?�q�q�?      �?      �?      �?              �?      �?              �?      �?              �?              �?        '!����?���n��?�������?�������?      �?                      �?�yCސ�?8�yC��?/�袋.�?F]t�E�?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ^Cy�5�?Cy�5��?              �?      �?        >����?|���?      �?              �?      �?�؉�؉�?;�;��?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�Y7�"��?L�Ϻ��?�������?�?�$I�$I�?n۶m۶�?F]t�E�?]t�E�?      �?                      �?              �?333333�?333333�?ZZZZZZ�?�������?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        /�袋.�?F]t�E�?333333�?�������?      �?      �?              �?      �?                      �?      �?              �?        �������?�������?���{��?�B!��?'vb'vb�?�;�;�?UUUUUU�?UUUUUU�?      �?                      �?333333�?333333�?<<<<<<�?�?      �?        ۶m۶m�?�$I�$I�?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �������?�������?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ,�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K녔h2h3h4hph<�h=Kub��������       f                     @>AU`�z�?�           8�@                                �J+@���H.�?�            �r@               
                    �?0B��D�?(            �M@               	                   �B@؇���X�?             ,@                               `f�)@$�q-�?
             *@       ������������������������       �                      @                                   ;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                  �)@��S�ۿ?            �F@                                   �? �q�q�?             8@        ������������������������       �                     �?                                   4@�nkK�?             7@                                  �2@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     1@                                �|�=@�����?             5@                                �|Y;@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@               O                    �?��Vk���?�             n@              $                    �?�E��
��?m            �c@                                    �?��.N"Ҭ?.            @Q@       ������������������������       �        "             K@                                   �?�r����?             .@        ������������������������       �                      @               #                   �E@8�Z$���?
             *@              "                   �7@�8��8��?	             (@                !                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        %       >                    �?�.�+��??            �U@        &       5                 м�J@����"�?             =@       '       *                 ��";@      �?             0@        (       )                     �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        +       ,                 ���<@8�Z$���?             *@        ������������������������       �                     @        -       4                    H@�<ݚ�?	             "@       .       3                    C@�q�q�?             @       /       2                 �|?@z�G�z�?             @       0       1                 ��2>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        6       7                   �8@��
ц��?
             *@        ������������������������       �                      @        8       =                   �H@���|���?             &@       9       <                 X�,@@�<ݚ�?             "@        :       ;                 Ȫ�c@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ?       @                 ��$:@�BbΊ�?'             M@        ������������������������       �        	             0@        A       B                    �?X�Cc�?             E@        ������������������������       �                     �?        C       N                     �?��]�T��?            �D@       D       E                   �;@�n_Y�K�?            �C@        ������������������������       �                     @        F       I                   �>@�t����?             A@        G       H                   @L@"pc�
�?	             &@       ������������������������       �                     "@        ������������������������       �                      @        J       K                   �B@�nkK�?             7@        ������������������������       �                     &@        L       M                 03�U@�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                      @        P       W                    �?ܻ�yX7�?2            @U@        Q       R                    �?r�q��?             8@        ������������������������       �                     (@        S       V                     �?�8��8��?             (@       T       U                   �4@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        X       _                    �?(��+�?$            �N@       Y       ^                     �?@��8��?             H@        Z       [                 ���^@�����H�?             "@       ������������������������       �                     @        \       ]                    )@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �C@        `       a                    :@��
ц��?	             *@        ������������������������       �                     @        b       e                 ��X@�<ݚ�?             "@       c       d                    0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        g       �                    �?,�+Ά1�?�            �y@        h       �                 �|�=@\�sե��?E            �\@       i       �                 03�:@X&$�E�?:            �X@       j       �                 ��$1@r�q��?8             X@       k       n                   �0@j���� �?2            @U@        l       m                    %@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        o       �                    �?��%��?-            �R@        p       w                    <@� �	��?             9@        q       v                   �6@      �?              @        r       s                 �{@�q�q�?             @        ������������������������       �                     �?        t       u                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        x       }                    �?j���� �?             1@        y       z                    �?r�q��?             @        ������������������������       �                     @        {       |                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ~                        �|Y=@�eP*L��?             &@        ������������������������       �                      @        �       �                 �?$'@�q�q�?             "@       �       �                 ���@؇���X�?             @        ������������������������       �                     @        �       �                   @@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?ڡR����?            �H@       �       �                 ���@\-��p�?             =@        ������������������������       �                      @        �       �                    �?�>����?             ;@       ������������������������       �                     9@        ������������������������       �                      @        �       �                 ��(@z�G�z�?             4@       �       �                  ��@      �?	             0@        ������������������������       �                     @        �       �                 �|Y=@�	j*D�?             *@        ������������������������       �                     �?        ������������������������       �      �?             (@        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     0@        �       �                    �?P�0�e��?�            �r@       �       �                 �T)D@�E���?�            `l@       �       �                 �?�@@�@+��?�            �k@       �       �                   �:@ d�=��?E            @\@       �       �                    �?�y��*�?#             M@        ������������������������       �                     @        �       �                 ���@ pƵHP�?             J@        �       �                 ���@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �F@        �       �                 ��L@ �Jj�G�?"            �K@        ������������������������       �                     =@        �       �                 �Yu@ ��WV�?             :@        �       �                    >@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        �       �                 @3�@��2(&�??            �[@        �       �                   �9@      �?             0@        ������������������������       �                      @        �       �                    �?և���X�?             ,@        ������������������������       �                     �?        �       �                   �=@�n_Y�K�?             *@        ������������������������       �                     �?        �       �                   �?@�q�q�?             (@        ������������������������       �                     �?        �       �                   �A@���|���?             &@        ������������������������       �      �?             @        ������������������������       �����X�?             @        �       �                 `�X!@��8��)�?7            �W@        �       �                   �0@ �q�q�?             H@        ������������������������       �                     �?        �       �                    <@`Ql�R�?            �G@        �       �                 pf� @�IєX�?
             1@        ������������������������       �                      @        �       �                   �:@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     >@        �       �                 �|=@*
;&���?             G@        �       �                   �2@ 7���B�?             ;@        �       �                 �y�+@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     9@        �       �                   �?@�����?             3@       �       �                 �|�=@��
ц��?             *@       �       �                    �?�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�;@      �?             @        ������������������������       �                      @        �       �                 �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    #@�G�5��?.            @Q@        �       �                 ���4@`՟�G��?             ?@        ������������������������       �                     &@        �       �                    �?R���Q�?             4@        ������������������������       �                      @        �       �                    �?      �?             (@       �       �                    @      �?              @        �       �                 `f�:@      �?             @        ������������������������       �                     �?        �       �                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 pf�C@      �?             @        �       �                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @�˹�m��?             C@       ������������������������       �                     ?@        �       �                    �?և���X�?             @       �       �                    @���Q��?             @       �       �                   �C@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������.���|�?ӣ���?�z�G��?���(\��?�A�I��?��}ylE�?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?              �?�������?�������?      �?                      �?      �?        �������?�?�������?UUUUUU�?      �?        �Mozӛ�?d!Y�B�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?        =��<���?�a�a�?�������?�������?      �?                      �?      �?        ��ƕ���?5�5��?��؉���?;�;��?ہ�v`��?�3J���?              �?�?�������?              �?;�;��?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �f��o�?�2)^ �?	�=����?�i��F�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?;�;��?      �?        9��8���?�q�q�?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �؉�؉�?�;�;�?      �?        F]t�E�?]t�E]�?�q�q�?9��8���?�������?333333�?              �?      �?                      �?      �?        �{a��?���=��?      �?        %I�$I��?�m۶m��?      �?        KԮD�J�?jW�v%j�?;�;��?ى�؉��?              �?�������?�������?F]t�E�?/�袋.�?              �?      �?        �Mozӛ�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?      �?              �?        ;ڼOq��?q�����?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�;�;�?�؉�؉�?              �?9��8���?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?        �����?6�&f�1�?�9E[�?�~]R��?;Cb�ΐ�?b�ΐ���?UUUUUU�?UUUUUU�?ZZZZZZ�?�������?F]t�E�?]t�E�?      �?                      �?}���g�?���L�?�Q����?)\���(�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?        ZZZZZZ�?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?                      �?����X�?����S��?�{a���?a����?      �?        h/�����?�Kh/��?              �?      �?        �������?�������?      �?      �?      �?        vb'vb'�?;�;��?              �?      �?      �?      �?                      �?      �?              �?        �u�)�Y�?�)�Y7��?��z��U�?`�(tSR�?������?;Ӹ�Qg�?���	��?x�!���?�4�rO#�?GX�i��?              �?'vb'vb�?;�;��?۶m۶m�?�$I�$I�?      �?                      �?      �?        k߰�k�?��)A��?      �?        O��N���?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��.���?t�E]t�?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?;�;��?ى�؉��?      �?        �������?�������?              �?]t�E]�?F]t�E�?      �?      �?�m۶m��?�$I�$I�?�Q�٨��?br1���?�������?UUUUUU�?              �?}g���Q�?W�+�ɕ?�?�?      �?        �q�q�?�q�q�?      �?                      �?      �?        ���,d!�?8��Moz�?	�%����?h/�����?      �?      �?              �?      �?              �?        Q^Cy��?^Cy�5�?�;�;�?�؉�؉�?ffffff�?333333�?              �?      �?                      �?      �?              �?      �?              �?      �?      �?      �?                      �?��v`��?�%~F��?�1�c��?�s�9��?              �?333333�?333333�?      �?              �?      �?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?      �?      �?                      �?      �?        ��P^Cy�?^Cy�5�?      �?        �$I�$I�?۶m۶m�?�������?333333�?      �?      �?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJf��'hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                 ��.@>AU`�z�?�           8�@              #                     @ d��0u�?�            �v@                                   �?      �?2             R@                                   �?      �?             8@        ������������������������       �                      @                                  �J@��2(&�?             6@                               `f�)@P���Q�?             4@        ������������������������       �                     "@        	                          �*@�C��2(�?             &@       
                           �?      �?              @                                 @<@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                  �)@      �?!             H@                                  5@HP�s��?             9@                                  �2@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     4@                                �|�<@�㙢�c�?             7@        ������������������������       �                     $@                                �|�=@�	j*D�?	             *@        ������������������������       �                      @               "                   �*@"pc�
�?             &@                                  @@      �?              @        ������������������������       �                      @                                   C@�q�q�?             @        ������������������������       �                     �?                !                   �F@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        $       3                 �ٝ@�q�q�?�             r@        %       &                 03�@��GEI_�?'            �N@        ������������������������       �                     :@        '       (                    �?(N:!���?            �A@        ������������������������       �                      @        )       *                   �4@�FVQ&�?            �@@        ������������������������       �                     �?        +       2                 �Y�@      �?             @@       ,       -                 ���@�}�+r��?             3@       ������������������������       �                     "@        .       /                 �|�:@ףp=
�?             $@        ������������������������       �                     @        0       1                 �|�=@؇���X�?             @       ������������������������       �r�q��?             @        ������������������������       �                     �?        ������������������������       �        	             *@        4       a                 @3�@�������?�            `l@        5       @                    �?p�ݯ��?J            �\@        6       7                 �|Y=@X��ʑ��?            �E@        ������������������������       �                     @        8       9                    �?�Gi����?            �B@        ������������������������       �                     ,@        :       ?                 X��A@�nkK�?             7@       ;       >                 ��(@���N8�?             5@       <       =                 ���@$�q-�?	             *@        ������������������������       �                     @        ������������������������       �r�q��?             @        ������������������������       �                      @        ������������������������       �                      @        A       X                 �?�@����O��?0            �Q@       B       W                 �Yu@&y�X���?*             M@       C       N                    �?<ݚ)�?             B@        D       M                 �|�;@�q�q�?	             (@       E       F                 ���@�z�G��?             $@        ������������������������       �                     @        G       L                 �&B@      �?             @       H       I                    4@      �?             @        ������������������������       �                      @        J       K                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        O       P                 �|�<@r�q��?             8@       ������������������������       �                     2@        Q       R                 ��@�q�q�?             @        ������������������������       �                     �?        S       T                 �|Y>@z�G�z�?             @        ������������������������       �                      @        U       V                 �&B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        Y       \                   �=@�θ�?             *@        Z       [                    8@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ]       ^                   �?@�����H�?             "@        ������������������������       �                     @        _       `                   �A@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        b       �                    �?4��Q���?J            @\@       c       d                   �*@���2j��?@            �Y@        ������������������������       �                      @        e       n                 ���"@�ڊ�e��?>             Y@       f       g                    �?$Q�q�?(            �O@        ������������������������       �                     @        h       m                 ��i @ 	��p�?&             M@       i       l                   �3@�ʈD��?            �E@        j       k                   �1@�q�q�?             @        ������������������������       �      �?              @        ������������������������       �      �?             @        ������������������������       �                    �B@        ������������������������       �                     .@        o       v                 03S#@$G$n��?            �B@        p       q                   �<@�z�G��?             $@       ������������������������       �                     @        r       s                 �|Y=@      �?             @        ������������������������       �                      @        t       u                 �|�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        w       �                    �?�>����?             ;@       x       y                 ��&@؇���X�?             ,@        ������������������������       �                     @        z       {                 ��*@      �?              @        ������������������������       �                     �?        |                        ���,@؇���X�?             @        }       ~                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        �       �                 @�+@���!pc�?
             &@        �       �                    <@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                 ��-@؇���X�?             @       ������������������������       �                     @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                     @R�����?�            �u@       �       �                   �D@:u��|2�?�            p@       �       �                    �?��R[s�?t            �e@       �       �                    @@uvI��?<            �X@        �       �                     �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        :            �W@        �       �                   �<@և���X�?8            @S@        �       �                 �̰f@l��
I��?             ;@       �       �                    $@�+e�X�?             9@        ������������������������       �                     @        �       �                    7@�q�q�?             2@        �       �                  DW@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 0��I@d}h���?	             ,@       �       �                     �?      �?             @       �       �                   �;@      �?             @        ������������������������       �                     �?        �       �                 `f�D@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ��$:@ �o_��?$             I@        ������������������������       �        	             0@        �       �                 �D A@j���� �?             A@        �       �                 ���<@X�Cc�?             ,@       �       �                    �?      �?              @       �       �                     �?      �?             @       �       �                 ��";@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 03k:@      �?             @        ������������������������       �                     �?        �       �                 �|�?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|?@r�q��?             @       ������������������������       �                     @        �       �                     �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     �?      �?             4@       �       �                 p�w@�E��ӭ�?             2@       �       �                 �|Y>@�r����?             .@        ������������������������       �                     "@        �       �                   @K@�q�q�?             @        ������������������������       �                     @        �       �                 ��n^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?H�U?B�?1            �T@        �       �                    �?      �?             8@        �       �                    J@8�Z$���?             *@        �       �                    �?�q�q�?             @       �       �                 �D\J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                     �?�C��2(�?             &@        ������������������������       �                     @        �       �                   �8@r�q��?             @        ������������������������       �                      @        �       �                    �?      �?             @       �       �                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?\-��p�?!             M@        �       �                    �?�}�+r��?	             3@       �       �                   �H@@4և���?             ,@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        �       �                   �R@:�&���?            �C@       �       �                   �J@$G$n��?            �B@       �       �                 �T!@@�q�q�?             8@       �       �                   �H@     ��?
             0@       �       �                     �?�8��8��?             (@        �       �                   �F@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                      @        �       �                    �?"Ae���?;            �W@        �       �                    @��6���?             E@        �       �                    @r�q��?             @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��Y7@b�2�tk�?             B@       �       �                 @3�/@      �?             0@        ������������������������       �                     @        �       �                 �|�;@���|���?
             &@        �       �                     @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    A@ףp=
�?             4@       ������������������������       �        	             1@        �       �                   @C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �                       �T�I@      �?             J@                              �̌5@�����?            �H@                                �?�q�q�?             ;@                               @;@�r����?	             .@                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@                                 0@�q�q�?             (@        ������������������������       �                     @        	      
                   �?      �?              @       ������������������������       �                     @                                 +@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                 �?���7�?             6@       ������������������������       �                     &@                                 @�C��2(�?             &@                                  @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?DDDDDD�?�������?      �?      �?      �?      �?              �?t�E]t�?��.���?�������?ffffff�?              �?F]t�E�?]t�E�?      �?      �?�������?�������?      �?                      �?              �?              �?      �?              �?      �?q=
ףp�?{�G�z�?333333�?�������?      �?                      �?      �?        �7��Mo�?d!Y�B�?      �?        vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?              �?        UUUUUU�?�������?�d����?;ڼOqɰ?      �?        |�W|�W�?�A�A�?              �?>����?|���?              �?      �?      �?�5��P�?(�����?      �?        �������?�������?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?              �?        �����?{��U���?^Cy�5�?Cy�5��?�}A_�?��}A�?              �?o0E>��?#�u�)��?              �?�Mozӛ�?d!Y�B�?��y��y�?�a�a�?�؉�؉�?;�;��?      �?        �������?UUUUUU�?      �?              �?         �
���?�]�����?��FX��?�i��F�?��8��8�?�8��8��?�������?�������?333333�?ffffff�?              �?      �?      �?      �?      �?      �?              �?      �?              �?      �?                      �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �؉�؉�?ى�؉��?      �?      �?              �?      �?        �q�q�?�q�q�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?����	�?x�!���?�������?�������?              �?��Q��?
ףp=
�?~��}���?AA�?      �?        ������?�{a���?A_���?�}A_з?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?              �?        к����?���L�?ffffff�?333333�?      �?              �?      �?              �?      �?      �?      �?                      �?�Kh/��?h/�����?۶m۶m�?�$I�$I�?      �?              �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        F]t�E�?t�E]t�?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�ҁr},�?��F�i�?�g�g�g�?4�3�3��?PuPu�?X|�W|��?9/���?�Cc}h��?      �?      �?      �?                      �?              �?�$I�$I�?۶m۶m�?h/�����?Lh/����?���Q��?R���Q�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?۶m۶m�?I�$I�$�?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        
ףp=
�?�Q����?      �?        �������?ZZZZZZ�?�m۶m��?%I�$I��?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?              �?      �?      �?              �?      �?              �?      �?�q�q�?r�q��?�������?�?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �D�JԮ�?�v%jW��?      �?      �?;�;��?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?F]t�E�?]t�E�?              �?UUUUUU�?�������?              �?      �?      �?      �?      �?              �?      �?                      �?a����?�{a���?�5��P�?(�����?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �A�A�?�o��o��?к����?���L�?UUUUUU�?�������?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?              �?                      �?      �?              �?                      �?�w6�;�?W�+���?b�a��?=��<���?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�8��8��?9��8���?      �?      �?              �?F]t�E�?]t�E]�?�������?�������?      �?                      �?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?^N��)x�?����X�?UUUUUU�?UUUUUU�?�������?�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?              �?      �?      �?      �?              �?      �?              �?      �?        �.�袋�?F]t�E�?      �?        ]t�E�?F]t�E�?      �?      �?      �?                      �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJy"rhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM1hjh))��}�(h,h/h0M1��h2h3h4hph<�h=Kub������       r                 `f�$@�s�ˈ.�?�           8�@                                ���@�����?�            �p@        ������������������������       �                     A@               #                    �?:�&���?�            @m@                                   �?�s��:��?             C@                                   �?�t����?             1@        ������������������������       �                     �?               	                 ���@      �?             0@        ������������������������       �                     �?        
                        �|�9@��S�ۿ?             .@        ������������������������       �                     @                                03@�8��8��?	             (@                                  �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                   3@����X�?             5@                                  �1@      �?             @        ������������������������       �                     �?                                P��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               "                 `��!@@�0�!��?             1@              !                 `�X!@���!pc�?             &@                                P�@z�G�z�?             $@                                  8@�q�q�?             @        ������������������������       �                     �?                                  �9@z�G�z�?             @        ������������������������       �                      @                                P��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        $       %                 ��@ �Cc}�?�            �h@        ������������������������       �                      @        &       K                 �?�@t�[ܝ�?�            @h@       '       J                    �?Xl���?L            �\@       (       1                 �Y�@ (��?K            @\@        )       *                   �5@      �?             0@        ������������������������       �                     �?        +       ,                 ���@��S�ۿ?
             .@        ������������������������       �                     @        -       .                 �|=@ףp=
�?             $@        ������������������������       �                     @        /       0                 �|�=@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        2       3                 ���@h�a��?@            @X@        ������������������������       �        
             1@        4       ?                 �?$@      �?6             T@        5       :                    �?�C��2(�?            �@@       6       7                 �|Y=@�����H�?             2@        ������������������������       �                     �?        8       9                 X��A@�IєX�?             1@       ������������������������       �$�q-�?	             *@        ������������������������       �                     @        ;       >                 �|Y>@��S�ۿ?	             .@       <       =                 �|�;@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        @       A                   �<@`�q�0ܴ?!            �G@       ������������������������       �                     =@        B       E                    �?�����H�?             2@        C       D                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        F       I                 �Yu@@4և���?             ,@        G       H                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             (@        ������������������������       �                     �?        L       M                ��k @R���Q�?5             T@        ������������������������       �                     �?        N       q                   @@@p#�����?4            �S@       O       ^                   �<@�� =[�?,             Q@       P       ]                 @�!@�t����?             A@       Q       X                   �3@���y4F�?             3@        R       U                   �1@և���X�?             @        S       T                   �0@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        V       W                 0S5 @      �?             @        ������������������������       �                      @        ������������������������       �                      @        Y       Z                 pf� @�8��8��?	             (@       ������������������������       �                     "@        [       \                    8@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     .@        _       b                 �|Y=@H�V�e��?             A@        `       a                 ���"@      �?             @       ������������������������       �                      @        ������������������������       �                      @        c       h                 �|�=@r�q��?             >@       d       e                 ��) @�����H�?
             2@       ������������������������       �                     .@        f       g                 pf� @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        i       n                   �?@      �?             (@        j       m                   �>@���Q��?             @       k       l                 �̌!@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        o       p                 ��I @؇���X�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                      @        ������������������������       �                     &@        s                         �D@��yƑ��?           �{@       t       �                 0�"K@
;&����?�            �u@       u       �                 ���C@����?�            pq@       v       �                    �?:��au��?�            �n@       w       �                 `f�)@�lO���?]             c@        x       y                    �?     ��?             @@        ������������������������       �                     @        z       �                    �?���>4��?             <@        {       |                 pF%@��S�ۿ?             .@       ������������������������       �                     &@        }       ~                     @      �?             @        ������������������������       �                      @               �                    +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    &@$�q-�?             *@       �       �                    5@�C��2(�?             &@        ������������������������       �      �?              @        ������������������������       �                     "@        ������������������������       �                      @        �       �                    �?�q�q�?I             ^@        �       �                   �;@      �?             F@        �       �                     @      �?
             ,@       �       �                   �9@r�q��?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?              @        �       �                   �-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     @�r����?             >@       ������������������������       �        
             ,@        �       �                 ��1@      �?	             0@       �       �                    �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �4@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                     �?�A+K&:�?,             S@        �       �                 ���<@��S���?	             .@        �       �                 `f&;@      �?             @       �       �                 �|�<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?���|���?             &@        ������������������������       �                      @        �       �                   �<@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �>@      �?              @       �       �                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?f>�cQ�?#            �N@        �       �                   �:@����X�?	             5@        ������������������������       �                     @        �       �                     @r�q��?             2@       ������������������������       �                     (@        �       �                 �|Y<@      �?             @        ������������������������       �                     �?        �       �                  �v6@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��,@��(\���?             D@        �       �                 �|�<@؇���X�?             5@       ������������������������       �                     (@        �       �                 �|�=@�q�q�?             "@        ������������������������       �                     �?        �       �                    @@      �?              @        ������������������������       �                      @        �       �                   @B@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     3@        �       �                     @$)}�~z�?<            �W@        �       �                   �;@�'�`d�?            �@@       �       �                   �6@���7�?             6@       ������������������������       �                     1@        �       �                    *@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `C@�eP*L��?             &@       �       �                   @A@�q�q�?             "@       �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�p����?'            �N@        �       �                 03�-@z�G�z�?	             .@        ������������������������       �                     �?        �       �                    -@؇���X�?             ,@        ������������������������       �                     �?        �       �                    �?$�q-�?             *@       ������������������������       �                     "@        �       �                    @      �?             @       �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @�I� �?             G@       �       �                    @�X����?             F@        �       �                    �?�t����?
             1@        ������������������������       �                     @        �       �                    @�n_Y�K�?	             *@       �       �                 ��|2@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�>����?             ;@        �       �                    +@؇���X�?	             ,@        ������������������������       �                     �?        �       �                    �?$�q-�?             *@        �       �                  ��6@z�G�z�?             @       �       �                   �=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             *@        �       �                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @r٣����?            �@@       �       �                    �?�q�q�?             8@        ������������������������       �                      @        ������������������������       �        	             0@        ������������������������       �                     "@        �       �                    �?r٣����?-            �P@       �       �                     @@4և���?             E@       ������������������������       �                    �C@        ������������������������       �                     @        �                          �?r�q��?             8@       �                       0wQ@�G��l��?             5@        �       �                      @؇���X�?             @       ������������������������       �                     @                                  >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �?X�Cc�?	             ,@                                �?�q�q�?             (@             
                p�w@���Q��?             @                               �8@      �?             @        ������������������������       �                      @              	                Ȫ�c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                              �̾w@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @              $                    �?����X�?9            �X@                                �?�BE����?%             O@        ������������������������       �                     *@              #                   �?ZՏ�m|�?            �H@             "                  �R@���y4F�?             C@             !                  @J@r�q��?             B@                              �5L@�q�q�?             2@                               @I@d}h���?             ,@                               �F@�8��8��?             (@                              03�C@r�q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                  G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                      @        ������������������������       �                     &@        %      &                `f�)@tk~X��?             B@        ������������������������       �                     @        '      ,                   �?��a�n`�?             ?@        (      +                  �.@      �?              @       )      *                    @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        -      0                  �*@���}<S�?             7@        .      /                  �F@z�G�z�?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     *@        �*       h�h))��}�(h,h/h0M1KK��h2h3h4hVh<�h=Kub��������������0Ȍ��?��o��?���-��?\�՘H�?      �?        �A�A�?�o��o��?�k(���?��k(��?�?<<<<<<�?              �?      �?      �?      �?        �?�������?              �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?      �?                      �?�m۶m��?�$I�$I�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ZZZZZZ�?�������?F]t�E�?t�E]t�?�������?�������?UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        %I�$I��?۶m۶m�?              �?-O"Ӱ��?���fy�?��>���?��Gp�?H���?x�!���?      �?      �?              �?�������?�?      �?        �������?�������?      �?        �������?UUUUUU�?�������?�������?      �?        �D�a�Y�?���Id�?      �?              �?      �?]t�E�?F]t�E�?�q�q�?�q�q�?              �?�?�?�؉�؉�?;�;��?      �?        �������?�?۶m۶m�?�$I�$I�?      �?                      �?      �?        ��F}g��?W�+�ɥ?      �?        �q�q�?�q�q�?      �?      �?              �?      �?        n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?              �?        333333�?333333�?              �?7a~W��?�#{���?�������?�������?<<<<<<�?�?6��P^C�?(������?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        iiiiii�?ZZZZZZ�?      �?      �?      �?                      �?�������?UUUUUU�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?333333�?�������?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?�������?�������?      �?              �?        a������?>����?�Mozӛ�?Y�B��?�[�f��?}Hw2��?!�M!�?�_��e��?��P^Cy�?�P^Cy�?      �?      �?              �?n۶m۶�?I�$I�$�?�?�������?              �?      �?      �?              �?      �?      �?              �?      �?        �؉�؉�?;�;��?]t�E�?F]t�E�?      �?      �?      �?              �?        �������?�������?      �?      �?      �?      �?UUUUUU�?�������?              �?      �?      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �?�������?              �?      �?      �?F]t�E�?]t�E�?      �?                      �?333333�?�������?      �?                      �?y�5���?�k(���?�������?�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        F]t�E�?]t�E]�?              �?�q�q�?r�q��?              �?      �?      �?�������?�������?      �?                      �?      �?        ��!XG�?�u�y���?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?      �?        �������?333333�?      �?                      �?�������?333333�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?        �l�w6��?����
�?'�l��&�?6�d�M6�?F]t�E�?�.�袋�?              �?�������?�������?      �?                      �?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?�������?333333�?              �?      �?              �?                      �?ާ�d��?C��6�S�?�������?�������?      �?        �$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?              �?      �?      �?      �?      �?              �?      �?                      �?Y�B���?Nozӛ��?�E]t��?]t�E]�?�������?�������?              �?ى�؉��?;�;��?r�q��?�q�q�?              �?      �?                      �?�Kh/��?h/�����?۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?�������?�������?      �?      �?      �?                      �?      �?              �?              �?              �?      �?      �?                      �?>���>�?|���?UUUUUU�?UUUUUU�?              �?      �?              �?        |���?>���>�?�$I�$I�?n۶m۶�?              �?      �?        UUUUUU�?UUUUUU�?��y��y�?1�0��?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?%I�$I��?�m۶m��?�������?�������?333333�?�������?      �?      �?      �?              �?      �?              �?      �?                      �?�$I�$I�?۶m۶m�?      �?                      �?      �?              �?        �m۶m��?�$I�$I�?)��RJ)�?���Zk��?              �?�>4և��?9/����?6��P^C�?(������?�������?UUUUUU�?UUUUUU�?UUUUUU�?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?                      �?      �?      �?      �?                      �?      �?                      �?      �?        r�q��?9��8���?      �?        �c�1��?�s�9��?      �?      �?333333�?�������?              �?      �?                      �?ӛ���7�?d!Y�B�?�������?�������?      �?      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�A�'hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       j                     @>AU`�z�?�           8�@               W                    �?����-�?�            �r@                                  �?��*��?�            �k@                                  �6@�ȉo(��?9            �V@                                   �?<���D�?            �@@        ������������������������       �                     @                                  �2@PN��T'�?             ;@                                  L@�8��8��?             8@       	                          �9@�nkK�?             7@        
                          �'@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     �?                                   ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        %             M@               *                   �@@RB)��.�?[             `@                                   �?���C��?*            �J@                                ���<@�q�q�?	             (@        ������������������������       �                     @                                  �9@      �?              @        ������������������������       �                     �?                                    �?և���X�?             @                               �|Y<@�q�q�?             @        ������������������������       �                     �?                                ��2>@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                )                     �?������?!            �D@       !       $                   �;@ףp=
�?             4@        "       #                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        %       (                   �>@�X�<ݺ?             2@        &       '                   @>@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             "@        ������������������������       �                     5@        +       2                    �?�w�"w��?1             S@        ,       1                     �?��
ц��?             *@       -       .                   �A@�eP*L��?             &@        ������������������������       �                     @        /       0                 м�J@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        3       T                   �J@���N8�?*            �O@       4       G                     �?p�v>��?             �G@       5       6                   @C@����"�?             =@        ������������������������       �                     @        7       B                   �G@�	j*D�?             :@       8       A                   �F@�t����?             1@       9       :                   @D@z�G�z�?             $@        ������������������������       �                     �?        ;       >                   �E@�<ݚ�?             "@        <       =                  x#J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ?       @                 ���K@r�q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        C       D                 ���E@�q�q�?             "@       ������������������������       �                     @        E       F                 ���W@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        H       K                   @A@r�q��?             2@        I       J                    1@�q�q�?             @        ������������������������       �      �?             @        ������������������������       �                      @        L       S                   �*@�8��8��?
             (@       M       N                   �'@r�q��?             @        ������������������������       �                     �?        O       R                   �F@z�G�z�?             @        P       Q                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        U       V                   �R@      �?
             0@       ������������������������       �        	             .@        ������������������������       �                     �?        X       _                    �?���y4F�?/             S@       Y       Z                    �? i���t�?             �H@       ������������������������       �                     ;@        [       \                 p"$X@�GN�z�?             6@       ������������������������       �                     (@        ]       ^                 Ъ�c@      �?             $@        ������������������������       �                     @        ������������������������       �                     @        `       g                    �?�5��?             ;@       a       d                     �?��
ц��?             *@       b       c                 �̾w@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        e       f                    *@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        h       i                   �3@����X�?             ,@       ������������������������       �                     $@        ������������������������       �                     @        k       z                    @Ԡ��	�?�            �y@        l       o                    �?�P�*�?             ?@        m       n                 pVE5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        p       s                    �?��>4և�?             <@       q       r                 @3�2@�n_Y�K�?             *@        ������������������������       �                      @        ������������������������       �                     @        t       u                 `f�:@���Q��?             .@        ������������������������       �                     @        v       y                    @���Q��?             $@       w       x                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        {       �                    �?r�q?�?�             x@        |       �                 �̌@ �.�6��?:             W@        }       ~                 ���@(;L]n�?             >@        ������������������������       �                     (@               �                 ��@�X�<ݺ?             2@        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                  ��8@f���M�?(             O@       �       �                    �?
;&����?             G@        �       �                 ��.@      �?
             0@       �       �                   �0@�q�q�?             @        �       �                    �?�q�q�?             @       �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                 ���4@�q�q�?             >@       �       �                 �|Y>@��}*_��?             ;@       �       �                    3@      �?             0@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 @3�@8�Z$���?
             *@        �       �                 �?�@      �?             @        ������������������������       �                     �?        �       �                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                   @B@�eP*L��?             &@       �       �                 03�1@      �?              @        ������������������������       �                     @        �       �                 03C3@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     0@        �                          �?,Ӕ��?�            @r@       �       �                    �?lE�ދ��?�            pq@        �       �                    �?�%^�?            �E@       �       �                   �6@R���Q�?             D@        �       �                 ��y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �0@��hJ,�?             A@       �       �                 ���@��a�n`�?             ?@        ������������������������       �                     (@        �       �                   @@�S����?
             3@       �       �                 �|=@���!pc�?             &@        ������������������������       �                      @        �       �                 �|�=@�q�q�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �                          �?8��%���?�            �m@       �       �                 �T)D@�����?�            �k@       �       �                    7@Dw�&��?�            �j@        �       �                 @3�@ ������?&            �O@       ������������������������       �                    �B@        �       �                 0S5 @ ��WV�?             :@        �       �                    1@r�q��?             @        ������������������������       �                     @        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     4@        �       �                   @@@�h�*$��?_             c@       �       �                   �>@H�ՠ&��?F             [@       �       �                 �?$@�C��2(�?B            �X@        �       �                    �?@�0�!��?             A@        �       �                 �|Y=@؇���X�?
             ,@        ������������������������       �                      @        ������������������������       �        	             (@        �       �                 P��@z�G�z�?             4@       �       �                 ���@      �?	             0@       �       �                   �8@      �?              @        �       �                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|�;@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        �       �                 03�6@P�2E��?,            @P@       �       �                    �?�]0��<�?)            �N@        ������������������������       �                     @        �       �                   �;@h㱪��?&            �K@        �       �                 pf� @�8��8��?             (@       ������������������������       �                     @        �       �                   �:@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|Y=@ qP��B�?            �E@        ������������������������       �        	             ,@        �       �                 ��) @XB���?             =@       ������������������������       �                     4@        �       �                 pf� @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|�:@      �?             @        ������������������������       �                      @        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �&B@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                 P�@      �?              @        ������������������������       �                     �?        �       �                   �?@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?`���i��?             F@        ������������������������       �                     �?        �       �                   @C@ qP��B�?            �E@        ������������������������       �                     5@        �       �                 @3�@���7�?             6@        �       �                   �C@�C��2(�?             &@        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     &@        �                          >@����X�?             @                                 ;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             ,@              
                   @�θ�?             *@             	                   #@      �?             (@                              83�@@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?��g�`�?��L���?־a���?� O	��?h�h��?�~��?|���?|���?              �?h/�����?&���^B�?UUUUUU�?UUUUUU�?d!Y�B�?�Mozӛ�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?S֔5eM�?���)k��?\�琚`�?"5�x+��?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?�������?333333�?              �?      �?              �?        p>�cp�?������?�������?�������?      �?      �?      �?                      �?��8��8�?�q�q�?�q�q�?�q�q�?      �?                      �?      �?              �?        ���k(�?��k(��?�;�;�?�؉�؉�?]t�E�?t�E]t�?              �?      �?      �?      �?                      �?      �?        �a�a�?��y��y�?ڨ�l�w�?L� &W�?	�=����?�i��F�?              �?vb'vb'�?;�;��?<<<<<<�?�?�������?�������?      �?        9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        UUUUUU�?UUUUUU�?              �?333333�?�������?      �?                      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?        �������?�������?      �?      �?      �?                      �?      �?              �?              �?      �?      �?                      �?(������?6��P^C�?����X�?/�����?              �?]t�E�?�袋.��?              �?      �?      �?      �?                      �?/�����?h/�����?�;�;�?�؉�؉�?۶m۶m�?�$I�$I�?      �?                      �?UUUUUU�?�������?              �?      �?        �$I�$I�?�m۶m��?              �?      �?        6�ɧ��?��l��	�?�Zk����?�RJ)���?UUUUUU�?UUUUUU�?              �?      �?        I�$I�$�?۶m۶m�?ى�؉��?;�;��?              �?      �?        �������?333333�?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUU��?�������?�B����?����7��?�?�������?              �?�q�q�?��8��8�?�$I�$I�?۶m۶m�?              �?      �?                      �?��RJ)��?��Zk���?Y�B��?�Mozӛ�?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?                      �?UUUUUU�?UUUUUU�?_B{	�%�?B{	�%��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?;�;��?;�;��?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ]t�E�?t�E]t�?      �?      �?              �?      �?      �?      �?                      �?      �?              �?              �?        �B�
*�?��իW��?�Q�ojT�?�ru��\�?�}A_��?�}A_�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?KKKKKK�?�������?�s�9��?�c�1Ƹ?      �?        (������?^Cy�5�?F]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?��V'�?A�IݗǶ?�Ϻ���?v�)�Y7�?����\��?��0�?��}��}�?AA�?      �?        O��N���?;�;��?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        y�5���?6��P^C�?������?{	�%���?]t�E�?F]t�E�?ZZZZZZ�?�������?۶m۶m�?�$I�$I�?              �?      �?        �������?�������?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?      �?        UUUUUU�?UUUUUU�?_�^��?z�z��?\2�h��?;ڼOqɠ?      �?        ־a���?��)A��?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?                      �?��}A�?�}A_З?      �?        GX�i���?�{a���?      �?        �q�q�?�q�q�?              �?      �?              �?      �?      �?              �?      �?              �?      �?        �q�q�?r�q��?      �?              �?      �?              �?۶m۶m�?�$I�$I�?              �?      �?        F]t�E�?F]t�E�?      �?        ��}A�?�}A_З?      �?        �.�袋�?F]t�E�?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?              �?        �$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?        ى�؉��?�؉�؉�?      �?      �?�������?333333�?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������       N                    �?�����?�           8�@                                    @�M���?�            �p@                                  �?$�q-�?V            �a@                                0Cd=@���}<S�?             G@                                  �C@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �B@        	                           @,���$�?:            @X@        
                        ��1V@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                    �?=QcG��?8            �W@        ������������������������       �                    �C@                                  @4@lGts��?!            �K@                                  B@      �?             @@       ������������������������       �                     4@                                  �C@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@                                   D@��<b���?             7@                                 �;@؇���X�?             5@                                   7@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                      @               /                 ��,#@H������?N            @^@                                   �?�<ݚ�?            �F@        ������������������������       �                     6@               .                    �?\X��t�?             7@               !                 ���@�\��N��?             3@        ������������������������       �                     �?        "       %                    8@X�<ݚ�?             2@        #       $                   �2@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        &       '                   �9@      �?	             (@        ������������������������       �                     @        (       )                 �Y5@�q�q�?             "@        ������������������������       �                     @        *       +                    ;@      �?             @        ������������������������       �                      @        ,       -                 ��� @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        0       7                    �?&:~�Q�?1             S@        1       4                 ��.@      �?             8@        2       3                 P��+@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        5       6                 X�,A@؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @        8       =                    @�θ�?"             J@        9       <                    �?؇���X�?             @       :       ;                 @3�2@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        >       C                    �?�r����?            �F@        ?       @                 �|�;@      �?             0@       ������������������������       �                     $@        A       B                    D@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        D       M                    @ 	��p�?             =@       E       L                   �>@�C��2(�?             6@       F       G                    4@���N8�?             5@        ������������������������       �                     $@        H       K                 @34@�C��2(�?	             &@        I       J                 ��/@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        O       \                    #@20��?%           �{@        P       Q                   �;@��X��?             <@        ������������������������       �        	             *@        R       S                    �?���Q��?	             .@        ������������������������       �                     �?        T       U                     @X�Cc�?             ,@        ������������������������       �                     @        V       W                 ��T?@ףp=
�?             $@        ������������������������       �                     @        X       Y                     @z�G�z�?             @        ������������������������       �                      @        Z       [                 ���A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ]       �                     �?��[���?           0z@        ^       �                   �J@l�Ӑ���?=            �U@       _       �                   �G@8�A�0��?.            �P@       `       �                   �E@�b��[��?'            �K@       a       b                 ��<:@~�4_�g�?              F@        ������������������������       �                     @        c       x                    �?      �?             C@        d       w                    �?���Q��?             4@       e       l                  Y>@p�ݯ��?             3@        f       g                 �|�;@      �?             @        ������������������������       �                     �?        h       k                 X�,@@�q�q�?             @       i       j                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        m       v                 �̾w@������?             .@       n       s                    �?d}h���?             ,@       o       p                 0�HU@r�q��?             (@       ������������������������       �                     @        q       r                 �|Y;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        t       u                 �nc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        y       �                    �?b�2�tk�?             2@       z       {                 �|�<@ҳ�wY;�?             1@        ������������������������       �                     @        |       }                   `@@և���X�?
             ,@        ������������������������       �                     @        ~       �                   @B@�q�q�?             "@              �                 �|Y>@؇���X�?             @        ������������������������       �                     @        �       �                   @K@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 ���E@���!pc�?             &@        ������������������������       �                     @        �       �                   �H@      �?             @        ������������������������       �                     �?        �       �                 (�`X@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?���N8�?             5@        ������������������������       �                     "@        �       �                    R@�8��8��?
             (@       ������������������������       �        	             &@        ������������������������       �                     �?        �       �                   @E@�+Ĺ+�?�            �t@       �       �                 0SE @l������?�            �r@       �       �                    �?$�Q�\�?i             e@       �       �                     @3��e��?g            �d@        ������������������������       �                     �?        �       �                   @@@��Lɿ��?f            �d@       �       �                   �>@p�"�0�?[            �b@       �       �                   @4@��ׄ��?U            `a@        �       �                   �3@r�q��?             B@       �       �                 �?�@$�q-�?             :@       ������������������������       �                     6@        �       �                   �2@      �?             @       �       �                    1@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���Q��?             $@        ������������������������       �                      @        �       �                 P�@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?b �57�?A            �Y@        �       �                   @9@r�q��?             (@        ������������������������       �                     �?        �       �                 ���@�C��2(�?             &@        ������������������������       �                      @        �       �                 �|=@�����H�?             "@        ������������������������       �                      @        �       �                 �|�=@؇���X�?             @       ������������������������       �r�q��?             @        ������������������������       �                     �?        �       �                    �?0�>���?:            �V@        �       �                 �|Y;@�nkK�?             7@        ������������������������       �                      @        �       �                  s�@���N8�?             5@        ������������������������       �                      @        �       �                 ��(@$�q-�?             *@       ������������������������       ��8��8��?             (@        ������������������������       �                     �?        �       �                 �|Y=@�IєX�?.             Q@       ������������������������       �                    �B@        �       �                 ��) @��� ��?             ?@       �       �                 �|�=@h�����?             <@       �       �                  sW@ 7���B�?             ;@        �       �                 pf�@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �?@      �?             $@        �       �                 pff@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 P�@և���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        ������������������������       �                     1@        ������������������������       �                      @        �       �                   �D@ �#�Ѵ�?Y             `@       �       �                   �7@ ��+,��?V            @_@       �       �                    �?H��2�?B            @W@        �       �                 �|�;@�r����?             .@        �       �                     @      �?             @        ������������������������       �                      @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�C��2(�?	             &@        ������������������������       �                     @        �       �                   `3@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �@@ ���J��?6            �S@       �       �                    &@����e��?-            �P@        �       �                   �3@ ��WV�?             :@        �       �                     @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     D@        �       �                     @�8��8��?	             (@       �       �                   �'@      �?              @        ������������������������       �                      @        �       �                   �A@r�q��?             @       �       �                    1@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @@        �       �                     @      �?             @       �       �                    4@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     A@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub������������������?��܍��?���>��?�>����?;�;��?�؉�؉�?d!Y�B�?ӛ���7�?�q�q�?r�q��?              �?      �?                      �?���fy�?�,O"Ӱ�?UUUUUU�?UUUUUU�?              �?      �?        AL� &W�?x6�;��?              �?�־a�?�<%�S��?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?��Moz��?��,d!�?�$I�$I�?۶m۶m�?333333�?ffffff�?              �?      �?                      �?      �?        �0�~�4�?�g���e�?�q�q�?9��8���?              �?��Moz��?!Y�B�?y�5���?�5��P�?              �?r�q��?�q�q�?UUUUUU�?�������?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?      �?      �?                      �?              �?�k(���?�k(����?      �?      �?ffffff�?333333�?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?        ى�؉��?�؉�؉�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ������?�{a���?]t�E�?F]t�E�?��y��y�?�a�a�?      �?        ]t�E�?F]t�E�?      �?      �?      �?                      �?      �?                      �?      �?        Χ�Q���?�`i��T�?%I�$I��?n۶m۶�?              �?333333�?�������?              �?%I�$I��?�m۶m��?              �?�������?�������?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        CF�T�?�ͅ�Xſ?�7[�~��?/�I���?颋.���?/�袋.�?� O	��?־a��?/�袋.�?��.���?      �?              �?      �?333333�?�������?^Cy�5�?Cy�5��?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?wwwwww�?�?I�$I�$�?۶m۶m�?�������?UUUUUU�?      �?        333333�?�������?              �?      �?              �?      �?              �?      �?                      �?              �?9��8���?�8��8��?�������?�������?              �?۶m۶m�?�$I�$I�?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?              �?      �?              �?        t�E]t�?F]t�E�?              �?      �?      �?              �?333333�?�������?      �?                      �?��y��y�?�a�a�?      �?        UUUUUU�?UUUUUU�?      �?                      �?(፦ί�?���ˊ��?+�3�=l�?��c.��?)ݾ�z��?�	j*D�?6�'���?S&���?      �?        �������?rY1P»?�PM�\"�?�y���?�Ke{��?��$D�?�������?UUUUUU�?�؉�؉�?;�;��?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?        333333�?�������?              �?      �?      �?      �?                      �?��VC��?�H%�e�?�������?UUUUUU�?              �?]t�E�?F]t�E�?      �?        �q�q�?�q�q�?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?        ��=��=�?�!�!�?�Mozӛ�?d!Y�B�?      �?        ��y��y�?�a�a�?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?        �?�?      �?        �{����?�B!��?�m۶m��?�$I�$I�?	�%����?h/�����?      �?      �?      �?                      �?      �?              �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?�������?�������?      �?              �?        �/����?�}A_Ч?`��"���?����Mb�?�~�駟�?X`��?�������?�?      �?      �?      �?              �?      �?      �?                      �?]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?��-��-�?�A�A�?�>����?|���?O��N���?;�;��?�q�q�?�q�q�?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?      �?      �?        �������?UUUUUU�?      �?      �?      �?      �?      �?              �?              �?              �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJJ��hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       z                     @�,�٧��?�           8�@                                  �1@Y(���?�            �s@        ������������������������       �                     ;@               s                   �M@      �?�             r@                                 �:@�?'>���?�            �p@                                   �?ҐϿ<��?"            �N@                                 �7@(;L]n�?             >@       ������������������������       �                     .@        	       
                     �?��S�ۿ?             .@        ������������������������       �                     $@                                  �+@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?f���M�?             ?@                                   �?     ��?             0@                                   �?��
ц��?             *@                                 �8@      �?             (@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                   4@�r����?	             .@                                 �2@"pc�
�?             &@        ������������������������       �                     @                                  �'@      �?              @       ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @               8                    �?      �?�            �i@               #                    �?��O���?0            @U@                                   �F@�8��8��?             8@       ������������������������       �                     2@        !       "                 83F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        $       7                    :@\#r��?"            �N@       %       .                   @4@b�h�d.�?            �A@       &       '                   �'@P���Q�?
             4@        ������������������������       �                     @        (       -                    -@@4և���?             ,@       )       *                   �B@�C��2(�?             &@       ������������������������       �                     "@        +       ,                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        /       6                    �?�q�q�?	             .@       0       1                     �?X�Cc�?             ,@        ������������������������       �                     @        2       3                   �;@�eP*L��?             &@        ������������������������       �                     @        4       5                    D@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     :@        9       d                  x#J@��p��?P            @^@       :       c                    �?��0{9�??            �W@       ;       b                  �>@r�q��?9             U@       <       O                 ��$:@��a�n`�?,             O@       =       J                   @D@�:�^���?            �F@       >       ?                   �)@�}�+r��?             C@        ������������������������       �                     3@        @       I                   @A@�KM�]�?             3@       A       H                    @@8�Z$���?
             *@       B       G                 ��,@�C��2(�?             &@       C       F                 �|�=@�����H�?             "@        D       E                 �|�<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        K       L                     �?����X�?             @        ������������������������       �                      @        M       N                   @F@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        P       a                     �?j���� �?             1@       Q       Z                    D@      �?             0@       R       S                 ��";@"pc�
�?	             &@        ������������������������       �                     @        T       U                 �ܵ<@����X�?             @        ������������������������       �                     �?        V       Y                 �|Y=@r�q��?             @        W       X                   @>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        [       \                    �?z�G�z�?             @        ������������������������       �                     �?        ]       `                 `f�;@      �?             @       ^       _                   @G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                     $@        e       p                    �?X�<ݚ�?             ;@       f       o                 �U�T@�\��N��?             3@       g       l                 03�M@����X�?	             ,@       h       k                   �C@      �?              @       i       j                    A@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        m       n                 Ј�Q@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        q       r                 @��v@      �?              @       ������������������������       �                     @        ������������������������       �                      @        t       y                    �?���}<S�?             7@       u       v                    �?؇���X�?	             ,@        ������������������������       �                     �?        w       x                   �R@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     "@        {       �                   �0@L K6R�?	           �x@        |       �                   �-@~h����?(             L@       }       �                    @�q�����?#             I@       ~                        @3�4@�û��|�?             7@        ������������������������       �        	             (@        �       �                    �?"pc�
�?
             &@        ������������������������       �                     @        �       �                    @����X�?             @        ������������������������       �                     @        �       �                 ��T?@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 `fV6@��}*_��?             ;@        �       �                 �&�)@�q�q�?             .@        ������������������������       �                     @        �       �                    �?�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �      �?              @        �       �                    �?�θ�?�             u@        �       �                    �?�D����?9             U@        �       �                    �?      �?             <@        �       �                 `�@1@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 03�:@�����?             5@       ������������������������       �                     3@        ������������������������       �                      @        �       �                    �?4և����?(             L@       �       �                 �|Y=@r�q��?#             H@        �       �                    <@���Q��?             $@       �       �                   �6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   `3@�}�+r��?             C@       �       �                    �?������?             B@       �       �                 ���@���N8�?             5@       ������������������������       �                     &@        �       �                   @@ףp=
�?             $@        �       �                 �|�=@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �2@      �?              @        ������������������������       �                      @        �       �                 ��.@r�q��?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �@�h1�
U�?�            �o@        ������������������������       �                     .@        �       �                    �?�t�9�?�            �m@        �       �                 ��,#@4�.�A�?(            �O@        �       �                  s@      �?             4@        ������������������������       �                     @        �       �                    �?X�Cc�?             ,@       �       �                 ��� @�eP*L��?	             &@       �       �                 P��@      �?             $@       �       �                    8@X�<ݚ�?             "@        ������������������������       �                     @        �       �                 �&B@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @1@�%^�?            �E@       �       �                 �|Y=@8�A�0��?             6@       �       �                    3@      �?
             0@        ������������������������       �                     �?        �       �                 pff0@z�G�z�?	             .@       �       �                   �:@$�q-�?             *@       ������������������������       �                     $@        �       �                   �&@�q�q�?             @        ������������������������       �                     �?        �       �                   �*@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��Y.@r�q��?             @        �       �                 ���*@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��p@@�����?             5@       �       �                    @"pc�
�?             &@       �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �                   �>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �9@h�V���?t             f@        �       �                 @3�@���N8�?(            �O@       ������������������������       �                    �@@        �       �                   �2@ףp=
�?             >@        �       �                 pf� @�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     5@        �                       �T�E@ ���x�?L            @\@       �                          �?,�T�6�?G             Z@       �                         @@@�+�$f��?B            �X@       �       �                 ��) @6YE�t�?-            �P@       �       �                   �@�*/�8V�?             �G@        �       �                   �?@����X�?	             ,@       �       �                 pf�@�C��2(�?             &@        ������������������������       �                     @        �       �                 �&B@؇���X�?             @       �       �                 �|�;@r�q��?             @        ������������������������       �                      @        �       �                 �|Y>@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@Pa�	�?            �@@       ������������������������       �                     2@        �       �                 �|�>@��S�ۿ?             .@       ������������������������       �                     (@        ������������������������       ��q�q�?             @                               �|�>@�d�����?             3@                             pf� @     ��?             0@        ������������������������       �                      @                                 (@d}h���?
             ,@             	                ���"@      �?              @                                <@z�G�z�?             @                                �:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        
                        �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                              @3�@      �?             @@                             �?�@��S�ۿ?             .@       ������������������������       �        	             *@        ������������������������       �      �?              @        ������������������������       �        
             1@        ������������������������       �                     @                                 �?X�<ݚ�?             "@                                ;@      �?              @        ������������������������       �                     @                              �|�>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������&��jq�?:�g *�?��8BF�?�)���\�?              �?      �?      �?�1�v��?��y#�?mާ�d�?������?�?�������?              �?�?�������?              �?�������?�������?      �?                      �?��RJ)��?��Zk���?      �?      �?�;�;�?�؉�؉�?      �?      �?      �?                      �?      �?                      �?�������?�?/�袋.�?F]t�E�?      �?              �?      �?333333�?�������?      �?              �?              �?      �?�?�������?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?XG��).�?��:��?_�_��?;��:���?�������?ffffff�?              �?�$I�$I�?n۶m۶�?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?�m۶m��?%I�$I��?              �?]t�E�?t�E]t�?      �?              �?      �?              �?      �?                      �?              �?fP*L��?j�V���?m�w6�;�?L� &W�?�������?UUUUUU�?�c�1��?�s�9��?}�'}�'�?l�l��?�5��P�?(�����?      �?        �k(���?(�����?;�;��?;�;��?]t�E�?F]t�E�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?      �?        �m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?        ZZZZZZ�?�������?      �?      �?F]t�E�?/�袋.�?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?�������?�������?      �?              �?      �?      �?      �?      �?                      �?      �?              �?              �?              �?        r�q��?�q�q�?�5��P�?y�5���?�$I�$I�?�m۶m��?      �?      �?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?ӛ���7�?d!Y�B�?۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?      �?                      �?      �?        �?��DO�?���@va�?�m۶m��?%I�$I��?�p=
ף�?���Q��?��,d!�?8��Moz�?              �?/�袋.�?F]t�E�?      �?        �m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?_B{	�%�?B{	�%��?UUUUUU�?UUUUUU�?              �?]t�E�?t�E]t�?      �?                      �?      �?        UUUUUU�?�������?              �?      �?      �?ى�؉��?�؉�؉�?�0�0�?z��y���?      �?      �?�m۶m��?�$I�$I�?      �?                      �?�a�a�?=��<���?              �?      �?        %I�$I��?n۶m۶�?�������?UUUUUU�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?�5��P�?(�����?�q�q�?�q�q�?��y��y�?�a�a�?      �?        �������?�������?      �?      �?UUUUUU�?UUUUUU�?      �?              �?              �?              �?      �?              �?      �?              �?      �?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?        �N���t�?��b�X,�?      �?        n�wp��?G" >���?�,˲,��?��i��i�?      �?      �?              �?�m۶m��?%I�$I��?]t�E�?t�E]t�?      �?      �?�q�q�?r�q��?              �?�������?�������?      �?                      �?      �?                      �?              �?�}A_��?�}A_�?颋.���?/�袋.�?      �?      �?              �?�������?�������?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?UUUUUU�?�������?      �?      �?              �?      �?                      �?=��<���?�a�a�?/�袋.�?F]t�E�?�q�q�?�q�q�?      �?        �������?�������?      �?                      �?      �?      �?      �?                      �?      �?        �袋.��?/�袋.�?��y��y�?�a�a�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        	�����?��	���?ى�؉��?;�;��?�Cc}h�?/�����?'�l��&�?e�M6�d�?r1����?m�w6�;�?�m۶m��?�$I�$I�?]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?              �?                      �?|���?|���?      �?        �������?�?      �?        UUUUUU�?UUUUUU�?Cy�5��?y�5���?      �?      �?              �?I�$I�$�?۶m۶m�?      �?      �?�������?�������?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?�������?�?      �?              �?      �?      �?              �?        r�q��?�q�q�?      �?      �?              �?�������?�������?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�U�uhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K兔h2h3h4hph<�h=Kub��������       B                    �?��t���?�           8�@                                    @���"͏�?�            0p@                                  �?=0�_�?]             c@                                 �;@Hm_!'1�?=            �X@                                    �?     ��?             @@       ������������������������       �        
             2@                                   �?X�Cc�?	             ,@        ������������������������       �                      @        	       
                   �'@�q�q�?             (@        ������������������������       �                     @                                  �7@      �?              @        ������������������������       �                     @        ������������������������       �                     @                                03�>@���7�?*            �P@                                  L@$�q-�?            �C@                               03[;@�}�+r��?             C@                                 �E@�?�|�?            �B@       ������������������������       �                     ;@                                  @G@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ;@        ������������������������       �                     �K@               A                    A@��U��?A            �Z@              6                    �?`՟�G��?9            @W@              #                   �@�%o��?,            �P@               "                 pff@�>����?             ;@                                 s@      �?              @       ������������������������       �                     @                !                 �|Y:@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     3@        $       /                    �?�Q����?             D@       %       ,                 �|�<@      �?             :@       &       '                   �0@�t����?             1@        ������������������������       �                     @        (       +                    3@$�q-�?	             *@        )       *                 `F�+@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        -       .                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        0       1                    @և���X�?	             ,@        ������������������������       �                     @        2       3                    �?���Q��?             $@        ������������������������       �                     @        4       5                 ���4@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        7       @                    @���B���?             :@       8       ;                    �?�J�4�?             9@        9       :                 �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        <       ?                 ��l4@�����?
             5@        =       >                 �|�:@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        ������������������������       �                     �?        ������������������������       �                     *@        C       P                    @C��wU�?           @|@        D       E                   �;@��H�}�?             9@        ������������������������       �                     "@        F       K                    �?     ��?	             0@        G       H                 �D,C@�q�q�?             "@        ������������������������       �                     @        I       J                      @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        L       M                    �?؇���X�?             @       ������������������������       �                     @        N       O                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Q       �                 ��$:@�������?           �z@       R       q                    �?l,��?�            `s@        S       b                 ��K.@����1�?/            @R@       T       U                     @P���Q�?&             N@        ������������������������       �                     @        V       Y                 �|Y=@�h����?#             L@        W       X                   �<@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        Z       [                    �?`Ql�R�?            �G@        ������������������������       �                     4@        \       a                 X��A@ 7���B�?             ;@       ]       ^                 ���@�nkK�?             7@        ������������������������       �                     (@        _       `                 ��(@�C��2(�?	             &@       ������������������������       �ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     @        c       d                 ��.@�	j*D�?	             *@        ������������������������       �                     �?        e       f                 ��$1@      �?             (@        ������������������������       �                     @        g       h                     @      �?              @        ������������������������       �                      @        i       n                    �?      �?             @       j       k                   �2@      �?             @        ������������������������       �                     �?        l       m                 �|�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        o       p                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        r       s                    )@x,����?�            �m@        ������������������������       �                     @        t       �                 �|�=@�X�<ݺ?�            @m@       u       �                   �4@X�.�d�?\            �a@        v       �                    �?�C��2(�?             F@       w       z                   �0@�ʈD��?            �E@        x       y                 �̌!@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        {       |                 �?�@�8��8��?             B@        ������������������������       �                     &@        }       ~                   �1@H%u��?             9@        ������������������������       �                      @               �                 @3�@�LQ�1	�?             7@        ������������������������       �                     �?        �       �                 ��Y @�C��2(�?             6@        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    &@�X�<ݺ?
             2@       �       �                     @ףp=
�?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|Y=@@uvI��?@            �X@       ������������������������       �        &            @P@        �       �                     @Pa�	�?            �@@        �       �                     �?      �?              @        ������������������������       �                     @        �       �                    @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     9@        �       �                     @���}<S�?;             W@        �       �                   �D@ ���J��?            �C@       ������������������������       �                     6@        �       �                   �*@�IєX�?             1@        �       �                    G@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     $@        �       �                 �?�@^�!~X�?             �J@        ������������������������       �                     3@        �       �                 ���'@H�V�e��?             A@       �       �                   �@@j���� �?             1@        �       �                 �̌!@����X�?             @       �       �                   �>@      �?             @        ������������������������       �                     �?        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 @3�@z�G�z�?             $@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     1@        �       �                 �\@z)�J'c�?G            @]@       �       �                    �?^����?@            @Z@        �       �                    <@���>4��?             <@        �       �                 pVAH@���!pc�?             &@        �       �                 ��A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �8@      �?              @        �       �                   �7@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 м�J@�t����?             1@       ������������������������       �                     "@        �       �                 м�M@      �?              @        ������������������������       �                     @        �       �                    I@���Q��?             @       �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 03k:@���!pc�?,            @S@        ������������������������       �                      @        �       �                    R@��{�?6�?+            �R@       �       �                    �?x�� ���?*            @R@       �       �                     @��U/��?             �L@       �       �                   �<@���3�E�?             J@        �       �                    8@���|���?             &@        ������������������������       �                     @        �       �                   �;@      �?              @        ������������������������       �                      @        �       �                 `f�D@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    K@� ��1�?            �D@       �       �                    �?r֛w���?             ?@        ������������������������       �                     �?        �       �                 `f�;@������?             >@        �       �                 X��B@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @K@z�G�z�?             9@       �       �                 �T!@@�����H�?	             2@        �       �                   @>@      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    C@և���X�?             @        �       �                 `f�N@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    ;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             0@        ������������������������       �                      @        ������������������������       �                     (@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������nԾ���?5"W��6�?*�Y7�"�?v�)�Y7�?p�pŪ?��S��S�?9/���?Y�Cc�?      �?      �?              �?�m۶m��?%I�$I��?              �?�������?�������?              �?      �?      �?      �?                      �?F]t�E�?�.�袋�?;�;��?�؉�؉�?(�����?�5��P�?к����?*�Y7�"�?              �?�������?�������?      �?                      �?      �?              �?                      �?              �?�[�琚�?tHM0���?�s�9��?�1�c��?\�՘H�?���[��?h/�����?�Kh/��?      �?      �?              �?      �?      �?              �?      �?                      �?ffffff�?�������?      �?      �?�������?�������?              �?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?        �q�q�?�q�q�?      �?                      �?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��؉���?ى�؉��?�z�G��?{�G�z�?      �?      �?              �?      �?        =��<���?�a�a�?333333�?�������?              �?      �?              �?                      �?      �?        KO-����?��JO-��?
ףp=
�?{�G�z�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        S_#Ot��?��r�.�?�M�4��?���/Y��?�Ν;w��?Ĉ#F��?ffffff�?�������?      �?        �$I�$I�?۶m۶m�?9��8���?�q�q�?      �?                      �?}g���Q�?W�+�ɕ?      �?        	�%����?h/�����?�Mozӛ�?d!Y�B�?      �?        ]t�E�?F]t�E�?�������?�������?      �?              �?        vb'vb'�?;�;��?              �?      �?      �?      �?              �?      �?      �?              �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        Y�>���?;�
_H�?              �?��8��8�?�q�q�?�ۥ����?�@�6�?]t�E�?F]t�E�?A_���?�}A_з?۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        )\���(�?���Q��?      �?        ��Moz��?Y�B��?              �?]t�E�?F]t�E�?      �?      �?              �?      �?        ��8��8�?�q�q�?�������?�������?      �?      �?      �?              �?              �?        �Cc}h��?9/���?      �?        |���?|���?      �?      �?      �?        �������?�������?      �?                      �?      �?        ӛ���7�?d!Y�B�?��-��-�?�A�A�?      �?        �?�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?        �}�	��?�	�[���?      �?        iiiiii�?ZZZZZZ�?�������?ZZZZZZ�?�$I�$I�?�m۶m��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?�������?�������?      �?      �?      �?              �?        7k�6k��?�)��)��?6Z�5Z��?�K��K��?I�$I�$�?n۶m۶�?t�E]t�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?              �?      �?                      �?�������?�������?      �?              �?      �?              �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        F]t�E�?t�E]t�?              �?�K~���?7�i�6�?Ĉ#F��?�ܹs���?Lg1��t�?g1��t�?O��N���?b'vb'v�?F]t�E�?]t�E]�?      �?              �?      �?              �?UUUUUU�?�������?              �?      �?        ������?������?���{��?�B!��?      �?        wwwwww�?�?�������?333333�?      �?                      �?�������?�������?�q�q�?�q�q�?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?              �?              �?        333333�?�������?              �?      �?              �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW��]hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       H                    �?e�L��?�           8�@                                    @��}� �?�            �o@                                  �?��S�ۿ?[            �b@                                 �*@�^'�ë�?:            @X@                                `f�)@ �o_��?             9@                                 �J@      �?
             0@       ������������������������       �        	             .@        ������������������������       �                     �?        	       
                    ;@�q�q�?             "@        ������������������������       �                     @                                  �A@      �?             @       ������������������������       �                     @        ������������������������       �                     @                                0Cd=@ �q�q�?,             R@                                  �H@H%u��?             9@                                 �;@P���Q�?             4@                                   �?z�G�z�?             @        ������������������������       �                      @                                  �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             .@                                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �G@        ������������������������       �        !            �J@               G                  ��8@��B����?C             Z@              (                 �̌@�K��&�?8            �U@               %                    �?d}h���?             <@                                �|Y8@�IєX�?             1@        ������������������������       �                     @        !       $                 ���@�8��8��?             (@        "       #                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        &       '                   �7@�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        )       D                    �?l��[B��?&             M@       *       7                   �9@��B����?"             J@       +       0                  �#@�q�q�?             >@        ,       /                    �?z�G�z�?	             .@       -       .                    �?؇���X�?             ,@        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     �?        1       4                    �?��S���?
             .@        2       3                 �[$@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        5       6                    @      �?             $@        ������������������������       �                     @        ������������������������       �                     @        8       C                   @B@�GN�z�?             6@       9       <                 �|�<@�KM�]�?             3@        :       ;                   �;@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        =       >                    �?      �?	             0@        ������������������������       �                     @        ?       B                   �@@�����H�?             "@       @       A                 ��1@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        E       F                    @r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        I       T                    @��/T8�?"           �|@        J       K                    �?j���� �?
             1@        ������������������������       �                     @        L       M                    �?      �?             ,@        ������������������������       �                     @        N       S                     @�z�G��?             $@       O       P                     @      �?             @        ������������������������       �                     �?        Q       R                 ��!>@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        U       �                    �?��#:���?           �{@        V       u                  �	U@������?6            �V@       W       d                 ��K.@�7�QJW�?/            �R@       X       [                   �5@�:�^���?            �F@        Y       Z                 �{@      �?             @        ������������������������       �                      @        ������������������������       �                      @        \       c                 �|�=@������?            �D@       ]       ^                 �|=@�>����?             ;@        ������������������������       �                     $@        _       `                 ���@�t����?
             1@        ������������������������       �                     @        a       b                   @@z�G�z�?             $@       ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     ,@        e       t                    �?�z�G��?             >@       f       q                     @��X��?             <@       g       l                  Y>@��<b���?             7@        h       k                 X��@@և���X�?             @       i       j                 �ܵ<@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        m       p                 �|Y<@      �?
             0@        n       o                   �8@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        r       s                   �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        v                           �?������?             .@       w       z                 X�,@@      �?             (@        x       y                 �|Y;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        {       |                 @�pX@�����H�?             "@        ������������������������       �                     @        }       ~                   @E@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     �? �<#�?�            �u@        �       �                  i?@θ	j*�?&             J@        �       �                   �G@r�q��?             8@       �       �                   @B@�	j*D�?             *@       �       �                    <@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                 �̌*@      �?              @        ������������������������       �                      @        �       �                 `fF<@      �?             @        �       �                 �|�?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    L@���|���?             &@        ������������������������       �                     @        �       �                    R@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?d}h���?             <@       �       �                    �?      �?             8@        ������������������������       �                     �?        �       �                 03�S@��+7��?             7@       �       �                 �|Y>@R���Q�?             4@        ������������������������       �                     @        �       �                    F@d}h���?
             ,@        �       �                   �C@      �?              @       �       �                 `f�K@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �T�I@@�z���?�            �r@       �       �                    @�5�s��?�             r@       �       �                   �2@�����?�            �q@        �       �                    �?r٣����?            �@@       �       �                     @�X����?
             6@        ������������������������       �                     @        �       �                 ��Y @     ��?             0@        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�C��2(�?	             &@       ������������������������       �                      @        �       �                    $@�q�q�?             @       �       �                 83�@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                  ��@���[s�?�            �o@        ������������������������       �                    �F@        �       �                    �?X��J��?�             j@        �       �                   `3@�KM�]�?             3@       �       �                 ��(@�X�<ݺ?             2@       ������������������������       �@4և���?             ,@        ������������������������       �                     @        ������������������������       �                     �?        �       �                     @x
�==Q�?y            �g@        �       �                   �@@��ϭ�*�?"             M@        ������������������������       �                     9@        �       �                    �?6YE�t�?            �@@       �       �                   �E@�חF�P�?             ?@       �       �                   @D@�d�����?
             3@       �       �                   @A@؇���X�?             ,@        �       �                    1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    4@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �        	             (@        ������������������������       �                      @        �       �                 �?$@�FVQ&�?W            �`@        �       �                 �|Y>@����X�?             @       �       �                 �|Y9@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?H�Swe�?R            @_@       �       �                 �?�@����&!�?N            @^@        ������������������������       �                     @@        �       �                 @3�@���M�?8            @V@        �       �                   �=@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                 pf!@Ћ����?3            �T@        ������������������������       �                    �@@        �       �                 `�X#@��<D�m�?            �H@       �       �                 ���"@�S����?             3@       �       �                 ���!@�C��2(�?	             &@       �       �                 �|Y<@      �?              @        �       �                   �:@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �<@      �?              @        ������������������������       �                     @        �       �                 �|Y=@���Q��?             @        ������������������������       �                     �?        �       �                 �|�=@      �?             @        ������������������������       �                      @        �       �                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     >@        ������������������������       �                     @        ������������������������       �                     @        �       �                    ;@      �?              @        ������������������������       �                      @        �       �                 p�O@�q�q�?             @        �       �                    >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������v�S(��?��X��?�@ �?��~����?�?�������?���Id�?=�L�v��?�Q����?
ףp=
�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?�������?���Q��?)\���(�?�������?ffffff�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?333333�?      �?                      �?              �?              �?ى�؉��?O��N���?���)k��?��)kʚ�?۶m۶m�?I�$I�$�?�?�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?]t�E�?t�E]t�?              �?      �?        ���=��?GX�i���?O��N���?ى�؉��?UUUUUU�?UUUUUU�?�������?�������?۶m۶m�?�$I�$I�?              �?      �?                      �?�?�������?333333�?�������?              �?      �?              �?      �?              �?      �?        ]t�E�?�袋.��?(�����?�k(���?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?�q�q�?�q�q�?�������?�������?              �?      �?                      �?      �?        �������?UUUUUU�?              �?      �?              �?        ���͉�?�������?ZZZZZZ�?�������?              �?      �?      �?      �?        333333�?ffffff�?      �?      �?              �?333333�?�������?              �?      �?                      �?k߰��?�S�<%��?wwwwww�?�?t�@�t�?0��b�/�?}�'}�'�?l�l��?      �?      �?      �?                      �?p>�cp�?������?�Kh/��?h/�����?      �?        <<<<<<�?�?      �?        �������?�������?333333�?�������?      �?              �?        ffffff�?333333�?n۶m۶�?%I�$I��?��,d!�?��Moz��?�$I�$I�?۶m۶m�?�������?333333�?      �?                      �?      �?              �?      �?333333�?�������?      �?                      �?      �?        �������?�������?      �?                      �?      �?        �?wwwwww�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���&��?�4��g�?�؉�؉�?�N��N��?UUUUUU�?UUUUUU�?vb'vb'�?;�;��?r�q��?�q�q�?              �?      �?      �?      �?              �?      �?      �?      �?      �?                      �?      �?      �?      �?                      �?      �?        F]t�E�?]t�E]�?              �?�������?�������?      �?                      �?I�$I�$�?۶m۶m�?      �?      �?      �?        zӛ����?Y�B��?333333�?333333�?      �?        I�$I�$�?۶m۶m�?      �?      �?�������?UUUUUU�?      �?                      �?              �?      �?                      �?      �?        ��y���?}0T�1�?�d�&Jv�?��DɮM�?�fӍo�?_�d���?>���>�?|���?�E]t��?]t�E]�?      �?              �?      �?              �?      �?        ]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        ���p8�?����x<�?      �?        !ղ��?m�Vi�_�?�k(���?(�����?��8��8�?�q�q�?n۶m۶�?�$I�$I�?      �?                      �?���~��?Ai�
��?����=�?|a���?      �?        '�l��&�?e�M6�d�?�Zk����?��RJ)��?Cy�5��?y�5���?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?333333�?      �?      �?      �?              �?              �?        >����?|���?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        X9��v�?�~j�t��?Sa���i�?���!pc�?      �?        ��^����?�E(B�?�$I�$I�?۶m۶m�?      �?                      �?ԮD�J��?��+Q��?      �?        ��S�r
�?և���X�?(������?^Cy�5�?]t�E�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?      �?        333333�?�������?              �?      �?      �?      �?              �?      �?              �?      �?              �?              �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJt�mUhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       x                 `�X.@<C�`��?�           8�@              1                    �? �n���?�            �v@               *                   @B@P����?3             S@                                  �?���!pc�?,            �P@                                   �?���|���?             &@                               �|Y:@      �?              @                                   @؇���X�?             @        ������������������������       �                     @        	       
                   �,@      �?             @        ������������������������       �                      @                                  �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                P��+@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               )                 �|�=@^(��I�?$            �K@                                  �?f.i��n�?            �F@                                   �?�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?                                  �@����e��?            �@@        ������������������������       �                     @                                `fV$@|��?���?             ;@                                   �?�	j*D�?             *@       ������������������������       �                     "@        ������������������������       �                     @               (                    �?����X�?	             ,@                               pF%@�q�q�?             (@        ������������������������       �                     @                #                     @      �?              @        !       "                    :@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        $       %                    �?      �?             @        ������������������������       �                      @        &       '                   �;@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        +       0                     @z�G�z�?             $@       ,       -                   �D@      �?             @        ������������������������       �                     �?        .       /                   �J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        2       3                    ,@<����?�            �q@        ������������������������       �                     @        4       A                   �:@H�te�?�            `q@        5       <                 �Y�@�h����?C             \@        6       7                 ���@@4և���?             ,@       ������������������������       �        	             &@        8       9                   �2@�q�q�?             @        ������������������������       �                     �?        :       ;                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        =       @                   �0@@uvI��?7            �X@        >       ?                 �̌!@z�G�z�?             @       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        4            @W@        B       M                     @h7�R�
�?l            �d@        C       D                   �)@����?�?            �F@       ������������������������       �                     9@        E       F                    �?P���Q�?             4@        ������������������������       �                     �?        G       H                   �C@�}�+r��?             3@        ������������������������       �                     "@        I       L                   �*@ףp=
�?             $@        J       K                    G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        N       O                 ���@����W1�?R            @^@        ������������������������       �                     5@        P       w                   �C@�:pΈ��?E             Y@       Q       h                 �|�=@��{H�?=            �U@       R       ]                 �?$@<���D�?-            �P@        S       \                 ��@�θ�?             :@       T       W                 �|Y=@z�G�z�?             9@        U       V                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        X       Y                    �?��2(&�?             6@        ������������������������       �      �?             @        Z       [                 ���@�X�<ݺ?             2@        ������������������������       �                     @        ������������������������       ��8��8��?             (@        ������������������������       �                     �?        ^       _                 ��) @P���Q�?             D@       ������������������������       �                     8@        `       c                   �;@      �?             0@        a       b                 �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        d       e                 �|Y=@@4և���?	             ,@        ������������������������       �                     @        f       g                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        i       v                 ��)"@����X�?             5@       j       k                 �&B@���y4F�?             3@        ������������������������       �                     @        l       s                   @@@������?             .@        m       r                 @3�@և���X�?             @       n       o                   �@���Q��?             @        ������������������������       �                     �?        p       q                 �?�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        t       u                   @C@      �?              @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     *@        y       �                     @��(@��?�            �u@       z       �                    �?��*��?�            @n@       {       �                    :@T(y2��?H            �]@        |       �                  ��9@      �?             4@        }       �                   �;@ףp=
�?             $@       ~                          �6@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �E@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?Pa�	�?:            �X@       ������������������������       �        /            @S@        �       �                    �?��2(&�?             6@        ������������������������       �                     @        �       �                    @�S����?	             3@        ������������������������       �                     @        ������������������������       �                     0@        �       �                 p�w@������?G            �^@       �       �                 `ff:@@��,*�?E            �]@        �       �                 �z� @���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        �       �                  �>@j�Je���?9            �X@        �       �                   @>@
j*D>�?             :@       �       �                   �<@�G�z��?             4@       �       �                   �J@j���� �?
             1@       �       �                    @@���|���?             &@       �       �                 ��";@և���X�?             @        �       �                 �|�<@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     �?�<ݚ�?)             R@       �       �                    &@t�7��?#             O@        ������������������������       �                     @        �       �                   @H@(2��R�?"            �M@       �       �                   �G@&^�)b�?            �E@       �       �                    �?r�q��?             E@       �       �                    �?r�q��?             B@        �       �                   �A@�����H�?             "@        �       �                 X�lA@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                  x#J@�+$�jP�?             ;@       �       �                 �|�<@�IєX�?	             1@        ������������������������       �                     �?        ������������������������       �                     0@        �       �                 `f�N@���Q��?             $@        �       �                 `f�K@�q�q�?             @       �       �                 `�iJ@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �>@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                    L@      �?             $@       �       �                    �?����X�?             @       �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   �>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?����0�?I             [@        �       �                    �?�eP*L��?              F@        �       �                    �?@4և���?
             ,@       ������������������������       �                     $@        �       �                    @      �?             @       �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?d��0u��?             >@        �       �                 ���4@�q�q�?	             (@       �       �                    �?z�G�z�?             $@       �       �                 �|�;@      �?              @        ������������������������       �                     �?        �       �                 03�1@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    @r�q��?             2@       �       �                 `f7@z�G�z�?
             .@        ������������������������       �                      @        �       �                 ��T?@$�q-�?	             *@       ������������������������       �                     @        �       �                 ��p@@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��.@     ��?)             P@        ������������������������       �                     @        �       �                    3@r�q��?'             N@        �       �                    �? �q�q�?             8@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        �       �                 �J/@      �?             B@        ������������������������       �                     @        �       �                 �y�/@8^s]e�?             =@        ������������������������       �                     @        �       �                    �?z�G�z�?             9@       �       �                    �?�t����?             1@        �       �                  �v6@      �?             @       �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    9@8�Z$���?
             *@        ������������������������       �                     @        �       �                    ;@z�G�z�?             $@        ������������������������       �                     �?        �       �                 �|�>@�����H�?             "@       ������������������������       �                     @        �       �                 �T)D@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������܍�W�?/�F�JP�?j����p�?W�Lt�<�?Q^Cy��?�P^Cy�?t�E]t�?F]t�E�?F]t�E�?]t�E]�?      �?      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        J��yJ�?�7�}���?�>�>��?�`�`�?UUUUUU�?UUUUUU�?              �?      �?        6�d�M6�?e�M6�d�?              �?	�%����?{	�%���?vb'vb'�?;�;��?      �?                      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?                      �?              �?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ���%N�?�X�0Ҏ�?              �?�_��?���1O�?۶m۶m�?�$I�$I�?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �Cc}h��?9/���?�������?�������?      �?      �?      �?              �?        rY1P��?o4u~�!�?��I��I�?l�l��?      �?        ffffff�?�������?      �?        �5��P�?(�����?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ��eP*L�?���|���?      �?        ��Q���?�Q����?���C���?/�I���?|���?|���?ى�؉��?�؉�؉�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?��.���?t�E]t�?      �?      �?��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?ffffff�?�������?      �?              �?      �?      �?      �?              �?      �?        n۶m۶�?�$I�$I�?      �?              �?      �?              �?      �?        �m۶m��?�$I�$I�?6��P^C�?(������?      �?        wwwwww�?�?�$I�$I�?۶m۶m�?�������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��+��+�?����?fP*L��?����!p�?�5�5�?�F��F��?      �?      �?�������?�������?�������?�������?              �?      �?                      �?�������?333333�?              �?      �?        |���?|���?              �?t�E]t�?��.���?              �?^Cy�5�?(������?      �?                      �?�v%jW��?��+Q��?�e�e�?�5�5�?��y��y�?�a�a�?              �?      �?        x9/���?����>�?;�;��?b'vb'v�?�������?�������?�������?ZZZZZZ�?F]t�E�?]t�E]�?�$I�$I�?۶m۶m�?�������?333333�?              �?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?9��8���?�q�q�?SJ)��R�?��Zk���?              �?=�"h8��?'u_[�?���/��?�}A_��?�������?UUUUUU�?�������?UUUUUU�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        /�����?B{	�%��?�?�?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?UUUUUU�?              �?      �?                      �?      �?              �?      �?�$I�$I�?�m۶m��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�Kh/���?Lh/����?]t�E�?t�E]t�?�$I�$I�?n۶m۶�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?DDDDDD�?wwwwww�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?                      �?      �?        �������?UUUUUU�?�������?�������?              �?�؉�؉�?;�;��?      �?        �������?UUUUUU�?              �?      �?              �?              �?      �?              �?�������?UUUUUU�?�������?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?      �?        |a���?	�=����?              �?�������?�������?�������?�������?      �?      �?      �?      �?              �?      �?                      �?;�;��?;�;��?      �?        �������?�������?              �?�q�q�?�q�q�?      �?              �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJc��hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       V                    �?ʡ�;S��?�           8�@               3                  �>@É`���?_            �d@                               ��i @�q�q�?3            @W@                                   �?@�0�!��?             A@        ������������������������       �                     �?               	                   �6@6YE�t�?            �@@                                ��y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        
                        �|�=@ 7���B�?             ;@                               �|=@�8��8��?	             (@        ������������������������       �                     @                                ���@      �?              @        ������������������������       �                     @                                  @@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     .@               (                    �?�Ƀ aA�?            �M@                                 P,@�����?             C@                                   �?�q�q�?             (@        ������������������������       �                     @                                pF�#@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               !                 ���<@8�Z$���?             :@                                  �;@      �?
             0@                                  �8@      �?              @       ������������������������       �                     @                                �0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        "       '                   b>@�z�G��?             $@       #       &                     �?      �?             @       $       %                 X��E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        )       .                 ���.@�ՙ/�?             5@        *       -                    �?�q�q�?             (@       +       ,                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        /       0                    �?�����H�?             "@       ������������������������       �                     @        1       2                      @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        4       I                 p"�X@���"͏�?,            �R@       5       D                    �?(L���?            �E@       6       C                   @O@      �?             D@       7       <                 0�FF@�˹�m��?             C@        8       9                 `f�A@�q�q�?             @        ������������������������       �                     @        :       ;                 X�lC@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        =       >                  �}S@      �?             @@       ������������������������       �                     2@        ?       B                   �8@@4և���?             ,@        @       A                 0wKT@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        E       F                    �?�q�q�?             @        ������������������������       �                     �?        G       H                 pV�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        J       S                   �F@���@M^�?             ?@       K       N                    �?      �?             8@       L       M                    �?8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        O       P                  "&d@���|���?             &@        ������������������������       �                     @        Q       R                   �?@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        T       U                 ���f@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        W       �                    �?��hJ,��?e            �@        X       q                     @�ucQ?-�?n            @e@       Y       n                    L@<����?;            �W@       Z       i                    6@�ƫ�%�?9            @V@        [       \                    �?PN��T'�?             ;@        ������������������������       �                     �?        ]       h                   @4@8�Z$���?             :@       ^       _                   �'@�nkK�?             7@        ������������������������       �                     $@        `       g                   �+@$�q-�?             *@        a       f                    D@r�q��?             @       b       e                    �?�q�q�?             @       c       d                    B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        j       k                 ���a@0�z��?�?+             O@       ������������������������       �        %            �J@        l       m                    !@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        o       p                 �TF@      �?             @        ������������������������       �                     @        ������������������������       �                     @        r       y                    �?l�;�	�?3            �R@        s       x                 X�,A@�r����?             .@       t       u                 �|�9@@4և���?             ,@        ������������������������       �                     �?        v       w                 ���@$�q-�?
             *@        ������������������������       �                     �?        ������������������������       �        	             (@        ������������������������       �                     �?        z       {                    ,@�z�G��?'             N@        ������������������������       �                     &@        |       }                    3@f�Sc��?             �H@        ������������������������       �                     @        ~       �                 ���5@f.i��n�?            �F@              �                 �|Y=@*;L]n�?             >@       �       �                   �4@�E��ӭ�?             2@        ������������������������       �                     @        �       �                    ;@�q�q�?             .@       �       �                   �9@�q�q�?	             (@       �       �                    �?�z�G��?             $@       �       �                    7@�<ݚ�?             "@       �       �                   �5@���Q��?             @        �       �                 ��y!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 `f!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   @B@�q�q�?             (@       �       �                 03�1@�����H�?             "@       ������������������������       �                     @        �       �                 03C3@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��p@@��S�ۿ?             .@        �       �                 pVm<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                     �?t�[|��?�            `w@        �       �                    �?����e��?-            �P@       �       �                   �B@�ՙ/�?*            �O@        �       �                 ��$:@     ��?             @@        ������������������������       �                     @        �       �                   �>@��}*_��?             ;@       �       �                 `fF<@�X����?             6@       �       �                 �|�?@j���� �?	             1@        ������������������������       �                      @        �       �                   �K@�q�q�?             .@       �       �                   @G@�θ�?             *@       �       �                    D@�q�q�?             "@        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|�<@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                  x#J@��a�n`�?             ?@        ������������������������       �                     (@        �       �                 `�iJ@p�ݯ��?             3@        ������������������������       �                      @        �       �                    A@�t����?             1@        �       �                 �|Y>@և���X�?             @       �       �                    <@���Q��?             @        �       �                    7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?ףp=
�?             $@        ������������������������       �                     �?        �       �                    H@�����H�?             "@       ������������������������       �                     @        �       �                 ���W@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��) @�q{�A,�?�            @s@        �       �                 ���@�FVQ&�?[            �`@        ������������������������       �                     8@        �       �                 ���@�>����?I             [@        ������������������������       �                      @        �       �                  ��@ �h�7W�?H            �Z@        ������������������������       �        	             3@        �       �                    �? 	��p�??            �U@        �       �                 �|Y=@d}h���?
             ,@        ������������������������       �                      @        �       �                 X��A@�8��8��?	             (@       ������������������������       �ףp=
�?             $@        ������������������������       �                      @        �       �                 ��L@���(-�?5            @R@        ������������������������       �                     $@        �       �                   �@���N8�?/            �O@        �       �                    >@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �?�@h�����?)             L@        ������������������������       �                     3@        �       �                   �2@@-�_ .�?            �B@        ������������������������       �                     �?        �       �                 @3�@������?             B@        �       �                   �A@r�q��?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     >@        �       �                 �G�?D��2(�?o             f@        ������������������������       �                     @        �       �                    @��Po�'�?m            �e@        �       �                     @X�Cc�?             ,@        ������������������������       �                     �?        �       �                    �?�	j*D�?
             *@        ������������������������       �                     @        �       �                 ���9@���Q��?             $@        ������������������������       �                     @        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                    @      �?             @       �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �9@p`q�q��?b            �c@        ������������������������       �        #            �J@        �                          $@�r����??            @Z@        �                         �?@��S���?	             .@       �       �                   �<@���|���?             &@        �       �                   �;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �                        �|�=@؇���X�?             @       �       �                 ��)"@      �?             @       �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                  @����\�?6            �V@                               @A@�:�]��?            �I@              
                   �?��s����?             5@             	                   1@���y4F�?             3@                               �@@�q�q�?             (@       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     >@                                 ;@$�q-�?            �C@        ������������������������       �                     �?                                 �?�}�+r��?             C@                                `3@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                              �T�E@Pa�	�?            �@@       ������������������������       �                     >@                                 >@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������N���I5�?d�~`l��?\��l���?ұ�I���?UUUUUU�?UUUUUU�?ZZZZZZ�?�������?              �?'�l��&�?e�M6�d�?UUUUUU�?UUUUUU�?      �?                      �?	�%����?h/�����?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        ~ylE�p�?'u_�?Q^Cy��?^Cy�5�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?;�;��?;�;��?      �?      �?      �?      �?      �?              �?      �?      �?                      �?      �?        ffffff�?333333�?      �?      �?      �?      �?              �?      �?                      �?      �?        �a�a�?�<��<��?�������?�������?�q�q�?r�q��?      �?                      �?      �?        �q�q�?�q�q�?              �?      �?      �?      �?                      �?*�Y7�"�?v�)�Y7�?w�qG��?⎸#��?      �?      �?^Cy�5�?��P^Cy�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?�$I�$I�?n۶m۶�?UUUUUU�?�������?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �c�1��?�s�9��?      �?      �?;�;��?;�;��?              �?      �?        F]t�E�?]t�E]�?              �?�������?�������?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?�������?�������?�������?666666�?�X�0Ҏ�?���%N�?�as�ì?��x�3�?h/�����?&���^B�?              �?;�;��?;�;��?d!Y�B�?�Mozӛ�?              �?;�;��?�؉�؉�?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?              �?      �?        �B!��?|���{�?              �?�q�q�?�q�q�?      �?                      �?      �?      �?      �?                      �?ƒ_,���?t�@�t�?�?�������?�$I�$I�?n۶m۶�?              �?;�;��?�؉�؉�?      �?                      �?      �?        ffffff�?333333�?      �?        ����>�?������?              �?�`�`�?�>�>��?""""""�?�������?�q�q�?r�q��?      �?        UUUUUU�?UUUUUU�?�������?�������?ffffff�?333333�?9��8���?�q�q�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?              �?                      �?              �?      �?        UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?      �?      �?      �?                      �?      �?        �������?�?�������?�������?      �?                      �?      �?        �ٓ|�?�S����?e�M6�d�?6�d�M6�?�<��<��?�a�a�?      �?      �?      �?        B{	�%��?_B{	�%�?]t�E]�?�E]t��?ZZZZZZ�?�������?      �?        UUUUUU�?UUUUUU�?�؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?333333�?�������?              �?      �?        �c�1��?�s�9��?      �?        ^Cy�5�?Cy�5��?              �?�������?�������?۶m۶m�?�$I�$I�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�������?�������?      �?        �q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �S{��?�g�'Ĺ?>����?|���?      �?        �Kh/��?h/�����?              �?��sHM0�?"5�x+��?      �?        ������?�{a���?I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?        ��իW��?�P�B�
�?      �?        ��y��y�?�a�a�?۶m۶m�?�$I�$I�?      �?                      �?�m۶m��?�$I�$I�?      �?        S�n0E�?к����?              �?�q�q�?�q�q�?�������?UUUUUU�?      �?              �?      �?      �?        �E]t��?�袋.��?              �?qG�w�?w�qG�?%I�$I��?�m۶m��?              �?vb'vb'�?;�;��?      �?        333333�?�������?              �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?      �?                      �?      �?        T:�g *�?^-n����?      �?        �������?�?�?�������?F]t�E�?]t�E]�?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?                      �?              �?      �?        .؂-؂�?�>�>�?}}}}}}�?�?z��y���?�a�a�?6��P^C�?(������?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?        �؉�؉�?;�;��?              �?�5��P�?(�����?�������?�������?      �?                      �?|���?|���?      �?        UUUUUU�?UUUUUU�?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg�$hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM!hjh))��}�(h,h/h0M!��h2h3h4hph<�h=Kub������       z                     @|��;;��?�           8�@               Y                 �5L@d�����?�            `u@              R                    �?JV��|�?�            �n@                                  �?(Q����?z            @i@                                   �?��Zy�?            �C@        ������������������������       �                     *@                                    �?8�Z$���?             :@              	                 �|�;@������?             .@        ������������������������       �                      @        
                           H@8�Z$���?
             *@                                  C@�<ݚ�?             "@                               ��2>@      �?              @                                ���<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@               %                    �?�����?b            `d@                                  �;@�����H�?            �F@                                  �6@������?             .@        ������������������������       �                     @                                  �9@      �?              @                                  �3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  �/@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                                   �7@(;L]n�?             >@       ������������������������       �                     2@        !       $                   �=@�8��8��?             (@       "       #                    D@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        &       5                 ��$:@p/3�d��?F            �]@       '       (                     �?г�wY;�?+             Q@        ������������������������       �                     @        )       ,                    5@�g�y��?(             O@        *       +                   �2@      �?              @        ������������������������       �                     @        ������������������������       �      �?              @        -       4                   �*@@3����?$             K@       .       /                   �'@������?             B@        ������������������������       �                     1@        0       1                    @@�}�+r��?             3@        ������������������������       �                     $@        2       3                   @B@�����H�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     2@        6       E                    B@�z�G��?             I@        7       D                   @@@�G��l��?             5@       8       9                    7@j���� �?
             1@        ������������������������       �                      @        :       A                 `f�D@��S���?	             .@       ;       >                 �|Y=@����X�?             @        <       =                   `@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ?       @                 `fF<@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        B       C                 �!�I@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        F       Q                    R@\-��p�?             =@       G       P                    @@ �Cc}�?             <@       H       O                   �<@     ��?	             0@       I       N                 `f�:@�r����?             .@       J       M                    J@8�Z$���?             *@        K       L                   @G@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        S       T                   �6@>��C��?            �E@        ������������������������       �                     7@        U       V                    �?      �?             4@        ������������������������       �                     @        W       X                    �?      �?             0@       ������������������������       �                     $@        ������������������������       �                     @        Z       c                    �?�п�Sr�?6            @X@       [       \                    �?@3����?!             K@       ������������������������       �                     H@        ]       ^                    �?r�q��?             @        ������������������������       �                     �?        _       `                 ���[@z�G�z�?             @        ������������������������       �                      @        a       b                    )@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        d       y                   �H@X��ʑ��?            �E@       e       t                 �|Y>@<=�,S��?            �A@       f       g                    &@�eP*L��?             6@        ������������������������       �                     @        h       s                     �?�t����?	             1@       i       r                    :@�q�q�?             .@       j       o                    �?X�<ݚ�?             "@       k       l                 0�HU@      �?             @        ������������������������       �                     �?        m       n                 �U�X@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        p       q                 �nc@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        u       v                 ЈT@$�q-�?             *@        ������������������������       �                     @        w       x                 03�U@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        {       �                    �?���� �?�            w@        |       �                  ��@r�p���?K            �\@        }       �                    �?�n`���?             ?@       ~       �                 X��B@ �Cc}�?             <@              �                    �?�>����?             ;@       �       �                    �?�X�<ݺ?             2@        ������������������������       �                      @        �       �                 �|Y8@      �?             0@        ������������������������       �                     @        �       �                 ���@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                  s@�����H�?             "@        ������������������������       �                     @        �       �                 �|Y:@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��Bu��?6             U@       �       �                  �#@�'�=z��?*            �P@        �       �                   �9@z�G�z�?
             4@       �       �                    �?      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        �       �                    A@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|Y=@�LQ�1	�?              G@       �       �                    @\X��t�?             7@        �       �                 ��*4@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             0@       �       �                    �?���Q��?             $@        ������������������������       �                      @        �       �                    4@      �?              @       �       �                 `F�+@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    .@�LQ�1	�?             7@        �       �                 ��*@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|�=@P���Q�?             4@       ������������������������       �                     .@        �       �                   �>@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��T?@r�q��?             2@        ������������������������       �                     "@        �       �                 ��p@@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �                       �T�I@ ̈́Q���?�            �o@       �       	                   �?�o��gn�?�             o@       �       �                    �?������?�            `j@        �       �                   �6@�������?             A@        �       �                 ��y@���|���?             &@        ������������������������       �                      @        �       �                    '@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|Y=@���}<S�?             7@        �       �                   �<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|Y?@�X�<ݺ?             2@       �       �                   @@�C��2(�?	             &@       �       �                 ���@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �0@(+���?s             f@        �       �                 pFD!@����X�?             @        �       �                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?p��@���?n            @e@        �       �                  ��@�IєX�?
             1@        ������������������������       �                      @        �       �                 X��A@�����H�?             "@       �       �                 ��(@      �?              @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �?�@Բ r��?d             c@       �       �                    7@P��BNֱ?4            �T@        ������������������������       �                     5@        �       �                   �8@Hn�.P��?'             O@        �       �                 �&b@؇���X�?             @        ������������������������       �                     @        �       �                 `fF@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���@h㱪��?#            �K@        ������������������������       �                     8@        �       �                   �?@`Jj��?             ?@       �       �                 �|�<@ 7���B�?             ;@        ������������������������       �                      @        �       �                 �|Y>@�}�+r��?             3@       �       �                  sW@��S�ۿ?             .@        ������������������������       �      �?              @        ������������������������       �        	             *@        ������������������������       �                     @        �       �                 �&B@      �?             @        ������������������������       �                      @        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                       �|Y>@(N:!���?0            �Q@       �       �                   �:@�>����?%             K@       �       �                 0S5 @(;L]n�?             >@        �       �                 @3�@r�q��?             @        ������������������������       �                     �?        �       �                   �3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     8@        �       �                   �;@      �?             8@        ������������������������       �                     �?        �       �                 ��) @���}<S�?             7@        ������������������������       �                     &@        �       �                 pf� @r�q��?	             (@        ������������������������       �                     �?        �                          (@�C��2(�?             &@       �                        �|Y=@؇���X�?             @       �       �                   �<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                              @3�@      �?             0@                                �A@z�G�z�?             @                               �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     &@        
                         $@�d�����?             C@                                 �?��.k���?
             1@                                �?��
ц��?             *@                                �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                 @؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                              `f�9@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                 3@�����?             5@        ������������������������       �                     &@                                 7@z�G�z�?             $@        ������������������������       �                     �?                                 �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                                 ;@z�G�z�?             @        ������������������������       �                     @                                  >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0M!KK��h2h3h4hVh<�h=Kub������������|d�_Z�?�7s@K�?�A|��?x�A|�?���D�?���v��?��be�F�?
L:5r�?� � �?\��[���?              �?;�;��?;�;��?wwwwww�?�?              �?;�;��?;�;��?9��8���?�q�q�?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?              �?        J� P��?l	��_a�?�q�q�?�q�q�?�?wwwwww�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?              �?      �?        �?�������?              �?UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?      �?                      �?����c�?~ylE�p�?�?�?      �?        ��{���?�B!��?      �?      �?      �?              �?      �?���Kh�?h/�����?�q�q�?�q�q�?      �?        �5��P�?(�����?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?              �?        ffffff�?333333�?��y��y�?1�0��?�������?ZZZZZZ�?      �?        �?�������?�$I�$I�?�m۶m��?      �?      �?      �?                      �?�������?�������?      �?                      �?      �?      �?      �?                      �?              �?a����?�{a���?%I�$I��?۶m۶m�?      �?      �?�������?�?;�;��?;�;��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?                      �?qG�w��?$�;��?              �?      �?      �?      �?              �?      �?              �?      �?        ����?��AG��?h/�����?���Kh�?              �?UUUUUU�?�������?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?��}A�?�}A_�?X|�W|��?�A�A�?t�E]t�?]t�E�?              �?�������?�������?UUUUUU�?UUUUUU�?�q�q�?r�q��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?              �?      �?              �?              �?        ;�;��?�؉�؉�?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?        jW�v%j�?,Q��+�?�%��~�?m5x�@�?�c�1��?�9�s��?۶m۶m�?%I�$I��?h/�����?�Kh/��?�q�q�?��8��8�?              �?      �?      �?              �?�������?�������?      �?                      �?�q�q�?�q�q�?              �?�������?�������?              �?      �?              �?              �?        z��y���?�0�0�?|���?|��|�?�������?�������?      �?      �?      �?                      �?      �?      �?              �?      �?        d!Y�B�?Nozӛ��?!Y�B�?��Moz��?�$I�$I�?۶m۶m�?              �?      �?              �?      �?333333�?�������?              �?      �?      �?      �?      �?              �?      �?              �?              �?        Y�B��?��Moz��?UUUUUU�?UUUUUU�?              �?      �?        �������?ffffff�?              �?�������?�������?      �?                      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �j�Z�V�?�T*�J��?rY1P��?�7�:���?�.~��?w*���?�������?�������?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?      �?                      �?ӛ���7�?d!Y�B�?�������?�������?      �?                      �?��8��8�?�q�q�?]t�E�?F]t�E�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?        �?�x�?�^o�?�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�?�?�?      �?        �q�q�?�q�q�?      �?      �?      �?      �?      �?              �?        ^�]��?�g�g�?��FS���?���ˊ��?      �?        t�9�s�?�c�1ƨ?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ־a���?��)A��?      �?        ���{��?�B!��?	�%����?h/�����?      �?        �5��P�?(�����?�������?�?      �?      �?      �?              �?              �?      �?      �?              �?      �?              �?      �?        |�W|�W�?�A�A�?�Kh/��?h/�����?�������?�?�������?UUUUUU�?      �?        �������?�������?              �?      �?              �?              �?      �?              �?ӛ���7�?d!Y�B�?      �?        �������?UUUUUU�?              �?]t�E�?F]t�E�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        Cy�5��?y�5���?�������?�?�؉�؉�?�;�;�?�������?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?      �?              �?      �?        =��<���?�a�a�?      �?        �������?�������?              �?�q�q�?�q�q�?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�>D5hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                  x#J@��ҴҰ�?�           8�@                                  @��߫~�?~           �@                                   �?     ��?             @@                                 �C@�C��2(�?             6@                               ��*4@���N8�?             5@       ������������������������       �                     &@               
                    �?ףp=
�?             $@              	                     @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                    @�z�G��?             $@                                    @���Q��?             @        ������������������������       �                      @                                pf�@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   @z�G�z�?             @        ������������������������       �                     @                                `f�:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               {                 Ь�#@��k��e�?j           �@               :                    �?����;�?�            pq@               !                   �7@&:~�Q�?,             S@                                    �?"pc�
�?             &@                                  �?ףp=
�?             $@       ������������������������       �                     @                                �{@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        "       9                 �|Y?@
��[��?%            @P@       #       *                    �?�����?             �L@        $       %                    �?R���Q�?             4@        ������������������������       �                     �?        &       )                 �|Y=@�KM�]�?
             3@        '       (                   @@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        +       ,                 �|Y=@�Gi����?            �B@        ������������������������       �                      @        -       4                    �?<=�,S��?            �A@        .       /                 ���@؇���X�?             ,@        ������������������������       �                     @        0       3                 03@"pc�
�?             &@       1       2                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        5       6                 ���@���N8�?             5@        ������������������������       �                     @        7       8                 ��(@�IєX�?	             1@       ������������������������       �      �?             0@        ������������������������       �                     �?        ������������������������       �                      @        ;       z                    �?ܷ��?��?�            `i@       <       M                    �?ܴD��?�            @i@        =       F                   �@����X�?             5@        >       E                 �&B@      �?             $@       ?       @                 pf�@r�q��?             @        ������������������������       �                     �?        A       B                    4@z�G�z�?             @        ������������������������       �                      @        C       D                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        G       H                   �9@�C��2(�?             &@       ������������������������       �                     @        I       J                 �?�@      �?             @        ������������������������       �                      @        K       L                 @3�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        N       O                     @�����D�?u            �f@        ������������������������       �        	             0@        P       ]                 �?�@d#,����?l            �d@       Q       R                 ��@h�����?9             U@        ������������������������       �                    �D@        S       X                 �?$@Du9iH��?            �E@        T       W                 �|Y>@z�G�z�?             $@        U       V                 �|�;@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        Y       Z                    ?@Pa�	�?            �@@       ������������������������       �                     ?@        [       \                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ^       c                   �3@�
��P�?3            @T@        _       b                 0S5 @����X�?	             ,@        `       a                   �1@      �?              @        ������������������������       �      �?             @        ������������������������       �      �?             @        ������������������������       �                     @        d       o                 �|�=@pH����?*            �P@       e       h                 ��) @=QcG��?            �G@       f       g                   �4@      �?             @@        ������������������������       �      �?              @        ������������������������       �                     >@        i       j                 pf� @�r����?	             .@        ������������������������       �                     �?        k       n                 @3�!@@4և���?             ,@        l       m                    8@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        p       w                 ��)"@z�G�z�?             4@       q       v                 @3�@�t����?
             1@        r       u                   �A@���Q��?             @       s       t                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     (@        x       y                   �?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        |       �                    �?d��0u��?�            �r@        }       �                   �0@���e���?P            �_@        ~                            @b�2�tk�?	             2@        ������������������������       �                     @        �       �                    �?d}h���?             ,@        �       �                   �,@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?���?��?G            @[@       �       �                   �H@4?,R��?-             R@       �       �                     @��IF�E�?)            �P@       �       �                   �6@`���i��?             F@       �       �                   �;@���7�?             6@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                    8@      �?             @        ������������������������       �                      @        �       �                   �/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �        	             6@        �       �                 ���1@���!pc�?             6@       �       �                   �D@@�0�!��?
             1@       �       �                 �|�=@      �?	             0@       �       �                  S�-@�<ݚ�?             "@        �       �                 �[$@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�7@���Q��?             @        ������������������������       �                      @        �       �                 �|Y>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    K@      �?             @       �       �                     �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     @��%��?            �B@        ������������������������       �                     $@        �       �                    @��}*_��?             ;@       �       �                    �?�n_Y�K�?             :@        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                   �>@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @C@D�n�3�?             3@       �       �                 ��p@@�n_Y�K�?             *@       �       �                 �|Y=@z�G�z�?             $@        ������������������������       �                     @        �       �                 @3k;@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                     �?����M�?k            �e@        �       �                   �B@��f/w�?%            �N@       �       �                 ��$:@P����?             C@        ������������������������       �                     @        �       �                   �J@h+�v:�?             A@       �       �                   �G@|��?���?             ;@       �       �                    �?�q�q�?             8@       �       �                   @E@�eP*L��?             6@       �       �                    �?�\��N��?             3@        �       �                   @@@      �?             $@       �       �                   �<@r�q��?             @        ������������������������       �                     @        �       �                  Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�<@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                 X�,@@      �?              @       �       �                 `fF<@և���X�?             @        ������������������������       �                      @        �       �                   �>@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     7@        �       �                 ��.@@4և���?F             \@       �       �                 ��K.@Ԫ2��?$            �L@       �       �                   @A@lGts��?#            �K@       �       �                     @�S����?             C@       �       �                    &@z�G�z�?             >@        ������������������������       ��q�q�?             @        �       �                    �?PN��T'�?             ;@        ������������������������       �                     @        �       �                 �|Y;@r�q��?             8@       ������������������������       �        	             0@        �       �                 �|�=@      �?              @        ������������������������       �                     @        �       �                    @@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                      @        ������������������������       �        "            �K@        �       �                    �?      �?B             Y@       �       �                    �?�g�y��?(             O@       ������������������������       �        "             J@        �       �                      @z�G�z�?             $@       �       �                    �?�����H�?             "@        ������������������������       �                      @        �       �                 Ъ�c@؇���X�?             @        �       �                 ���[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �                         �E@\�Uo��?             C@       �                       �|Y>@�LQ�1	�?             7@       �                       �̰f@�n_Y�K�?             *@       �       �                   �1@�eP*L��?             &@        ������������������������       �                     @        �       �                     @      �?              @       �       �                   �9@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �        	             .@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub��������������(�TL�?���Vg�?���q�O�?����`�?      �?      �?F]t�E�?]t�E�?�a�a�?��y��y�?              �?�������?�������?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?        333333�?ffffff�?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?      �?              �?      �?        ��-�D�?����v�?�駟~�?X`��?�k(���?�k(����?F]t�E�?/�袋.�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        7r#7r#�?�����?Q^Cy��?^Cy�5�?333333�?333333�?              �?�k(���?(�����?      �?      �?      �?                      �?      �?        o0E>��?#�u�)��?              �?�A�A�?X|�W|��?�$I�$I�?۶m۶m�?              �?F]t�E�?/�袋.�?      �?      �?              �?      �?                      �?��y��y�?�a�a�?      �?        �?�?      �?      �?      �?              �?        ��=���?a���{�?�(0���?z��~�X�?�m۶m��?�$I�$I�?      �?      �?�������?UUUUUU�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?]t�E�?F]t�E�?      �?              �?      �?      �?              �?      �?              �?      �?        x�Y]��?>)7ͳ?      �?        I����H�?��[���?�m۶m��?�$I�$I�?      �?        qG�w��?w�qGܱ?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        |���?|���?      �?              �?      �?              �?      �?        ������?��ӭ�a�?�m۶m��?�$I�$I�?      �?      �?      �?      �?      �?      �?      �?        �1���?z�rv��?x6�;��?AL� &W�?      �?      �?      �?      �?      �?        �������?�?              �?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?      �?                      �?      �?        �������?�������?<<<<<<�?�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?                      �?DDDDDD�?wwwwww�?�d2�L&�?��f��l�?�8��8��?9��8���?              �?I�$I�$�?۶m۶m�?�������?333333�?              �?      �?              �?        N��ش�?-�M���?r�q��?�8��8��?'�l��&�?�l��&��?F]t�E�?F]t�E�?F]t�E�?�.�袋�?�������?�������?              �?      �?      �?              �?      �?      �?              �?      �?                      �?              �?t�E]t�?F]t�E�?�������?ZZZZZZ�?      �?      �?�q�q�?9��8���?      �?      �?              �?      �?                      �?              �?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?333333�?�������?      �?                      �?              �?}���g�?���L�?              �?_B{	�%�?B{	�%��?;�;��?ى�؉��?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?                      �?l(�����?(������?ى�؉��?;�;��?�������?�������?              �?�������?333333�?      �?                      �?      �?              �?              �?        (�j��?�6��<�?XG��).�?��!XG�?�P^Cy�?Q^Cy��?      �?        �������?xxxxxx�?{	�%���?	�%����?�������?�������?t�E]t�?]t�E�?�5��P�?y�5���?      �?      �?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?�q�q�?r�q��?              �?      �?      �?�$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?                      �?      �?              �?                      �?      �?              �?        n۶m۶�?�$I�$I�?$���>��?p�}��?�<%�S��?�־a�?(������?^Cy�5�?�������?�������?UUUUUU�?UUUUUU�?&���^B�?h/�����?      �?        �������?UUUUUU�?      �?              �?      �?              �?�������?�������?      �?              �?      �?      �?              �?                      �?      �?              �?      �?�B!��?��{���?              �?�������?�������?�q�q�?�q�q�?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �5��P^�?6��P^C�?d!Y�B�?Nozӛ��?;�;��?ى�؉��?t�E]t�?]t�E�?              �?      �?      �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���&hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       t                     @"��p�?�           8�@               k                    �?�h��?�             t@                                  �?�D�.1��?�            �q@                                  @L@�|1)�?G            �Z@                                  �?�q�q�?B             X@        ������������������������       �                     >@                                  �;@����e��?.            �P@               	                   �:@ 7���B�?             ;@       ������������������������       �                     9@        
                          �/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �C@                                  �L@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @               *                    �?���~X��?n            �f@               )                    I@r�qG�?             H@              &                    �?��Zy�?            �C@                                 @@@`՟�G��?             ?@                               ���<@      �?             4@        ������������������������       �                     $@                                �U�X@      �?             $@                               �|�;@r�q��?             @        ������������������������       �                     @                                03SA@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  �A@"pc�
�?             &@        ������������������������       �                     @                %                     �?���Q��?             @       !       "                   �A@      �?             @        ������������������������       �                      @        #       $                   @E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        '       (                 �̾w@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        +       ,                    #@���\�?T            �`@        ������������������������       �                     @        -       j                   �R@�nN@��?P            �_@       .       C                 ��D:@K�|%��?O            @_@       /       B                   �*@D��*�4�?*            @Q@       0       A                   @B@4��?�?!             J@       1       @                   �@@$G$n��?            �B@       2       ;                 `fF)@�#-���?            �A@       3       4                    @���7�?             6@        ������������������������       �                     @        5       :                    �?      �?             0@       6       9                    5@@4և���?
             ,@        7       8                   �2@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                      @        <       =                 �|�<@8�Z$���?             *@       ������������������������       �                     $@        >       ?                 �|�=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             .@        ������������������������       �        	             1@        D       i                    �?Dc}h��?%             L@       E       h                     �?�q�q�?!            �I@       F       a                   �G@�w��#��?              I@       G       R                   �>@0,Tg��?             E@        H       Q                 `f�<@�z�G��?             $@       I       J                 03k:@      �?              @        ������������������������       �                     �?        K       P                   �C@և���X�?             @       L       O                 �|�?@      �?             @       M       N                 �|�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                      @        S       X                 `fFJ@      �?             @@       T       W                 �|�<@ �q�q�?             8@        U       V                 `f�D@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             3@        Y       Z                    <@      �?              @        ������������������������       �                     �?        [       \                 �|Y>@����X�?             @        ������������������������       �                     @        ]       ^                 `f�K@      �?             @        ������������������������       �                     �?        _       `                    E@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        b       g                 ���T@      �?              @       c       f                    @@�q�q�?             @       d       e                    L@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        l       m                    @؇���X�?            �A@        ������������������������       �                      @        n       s                    B@�C��2(�?            �@@       o       r                    �?�g�y��?             ?@        p       q                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                      @        u       �                 �ٝ@;��t��?�            Px@        v       w                 ���@�8��8��?%             N@        ������������������������       �                     :@        x       y                    �?��hJ,�?             A@        ������������������������       �                      @        z       {                 ��@     ��?             @@        ������������������������       �                     �?        |       �                    �?`Jj��?             ?@       }       �                    �? 	��p�?             =@       ~       �                 ���@      �?
             0@              �                 �|�9@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 �|=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     *@        ������������������������       �                      @        �       �                    �?������?�            �t@        �       �                    �?�G�z��?3             T@        �       �                 ���@<���D�?            �@@        ������������������������       �                     �?        �       �                    �?     ��?             @@        �       �                    �?�q�q�?             "@       �       �                 �|�5@      �?              @       �       �                    @r�q��?             @        ������������������������       �                     @        �       �                 ��|*@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        �       �                 03s@��0{9�?            �G@        �       �                 �|Y=@���}<S�?             7@        ������������������������       �                      @        ������������������������       �                     5@        �       �                 �-!@�q�q�?             8@        ������������������������       �                     @        �       �                 �|Y<@�����?             5@        ������������������������       �                     (@        �       �                   `3@�<ݚ�?             "@       �       �                    �?؇���X�?             @       ������������������������       �                     @        �       �                 X�lA@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�4@*%�5P�?�             o@       �       �                    �?�:,&�e�?            �h@       �       �                   �@     ��?q             f@        �       �                    �?��V#�?            �E@        �       �                 �|�;@�t����?             1@       �       �                 pf�@z�G�z�?             .@        ������������������������       �                     @        �       �                 �&B@�z�G��?             $@        �       �                    4@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                 P�N@$�q-�?             :@       �       �                 �?$@P���Q�?             4@       �       �                 ��@�8��8��?	             (@        ������������������������       �                     @        �       �                 �|�;@؇���X�?             @        ������������������������       �                     @        �       �                 �|Y>@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        �       �                    >@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �?�@؇���X�?Y            �`@        ������������������������       �                     =@        �       �                    �?B�����?F             Z@        �       �                   �9@�z�G��?             4@       �       �                 ��&@�8��8��?	             (@       ������������������������       �                     $@        �       �                    '@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �A@      �?              @       �       �                 �|�;@r�q��?             @        ������������������������       �                      @        �       �                 pf�'@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 @3�@0,Tg��?6             U@        �       �                    :@�eP*L��?             &@        ������������������������       �                     @        �       �                   �A@����X�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                 `�X#@L������?0            @R@       �       �                    3@\-��p�?'             M@        �       �                   �1@�eP*L��?             &@       �       �                 pf� @�q�q�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���"@=QcG��?!            �G@       �       �                 @Q!@P�Lt�<�?             C@       ������������������������       �                     7@        �       �                    9@��S�ۿ?             .@        ������������������������       �                      @        �       �                    <@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �<@�<ݚ�?             "@        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�=@z�G�z�?             @        ������������������������       �                      @        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             .@        �       �                    �?��<b���?             7@       �       �                    �?�t����?             1@       �       �                   �;@�θ�?             *@       ������������������������       �                     @        �       �                 `fv1@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    &@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �                       �T�I@ףp=
�?             I@       �                         @C@P���Q�?             D@       �                         �B@@4և���?             <@       �                          @ 7���B�?             ;@        �                          �?ףp=
�?             $@                               ��T?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             1@        ������������������������       �                     �?        ������������������������       �                     (@                              �|�>@�z�G��?             $@             	                   �?      �?              @        ������������������������       �                     @        
                         ;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������J54v��?l�����?�.>9�?��h�`��?�9a��?cOy���?"5�x+��?W�9�&�?UUUUUU�?�������?              �?|���?�>����?h/�����?	�%����?              �?      �?      �?              �?      �?                      �?�������?�������?      �?                      �?�[#�˰�?"H��h��?�������?�������?� � �?\��[���?�1�c��?�s�9��?      �?      �?      �?              �?      �?UUUUUU�?�������?              �?      �?      �?              �?      �?              �?        F]t�E�?/�袋.�?              �?�������?333333�?      �?      �?              �?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?      �?        ��2.��?���7G��?              �?��(��(�?�u]�u]�?��|?5^�?�I+��?ہ�v`��?)�3J���?�N��N��?ى�؉��?к����?���L�?�A�A�?_�_�?�.�袋�?F]t�E�?      �?              �?      �?n۶m۶�?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?        ;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?��Q��?��(\���?�y��y��?1�0��?333333�?ffffff�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?�������?UUUUUU�?�������?�������?              �?      �?              �?              �?      �?              �?�m۶m��?�$I�$I�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?                      �?      �?              �?                      �?�$I�$I�?۶m۶m�?      �?        F]t�E�?]t�E�?�B!��?��{���?�q�q�?�q�q�?              �?      �?                      �?      �?        qD��C�?;�����?UUUUUU�?UUUUUU�?      �?        KKKKKK�?�������?              �?      �?      �?              �?���{��?�B!��?������?�{a���?      �?      �?]t�E�?F]t�E�?              �?      �?        �������?�������?      �?              �?      �?      �?              �?        %P�[:�?�_]H���?�������?�������?|���?|���?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?m�w6�;�?L� &W�?ӛ���7�?d!Y�B�?              �?      �?        UUUUUU�?�������?              �?=��<���?�a�a�?      �?        9��8���?�q�q�?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?      �?              �?      �?        ���[���?�������?��F���?~r!�f�?      �?      �?eMYS֔�?6eMYS��?�������?�������?�������?�������?              �?333333�?ffffff�?      �?      �?      �?                      �?              �?      �?        �؉�؉�?;�;��?ffffff�?�������?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?      �?              �?        �������?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?      �?        vb'vb'�?'vb'vb�?ffffff�?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        �0�0�?�<��<��?t�E]t�?]t�E�?      �?        �$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?�Ǐ?~�?����?a����?�{a���?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?x6�;��?AL� &W�?���k(�?(�����?      �?        �������?�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ��Moz��?��,d!�?�������?�������?�؉�؉�?ى�؉��?              �?      �?      �?      �?                      �?      �?      �?              �?      �?                      �?�������?�������?ffffff�?�������?n۶m۶�?�$I�$I�?	�%����?h/�����?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?      �?        ffffff�?333333�?      �?      �?      �?        �������?�������?              �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�EhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       d                    �?>AU`�z�?�           8�@               ]                 ���Q@�.�~��?�            �p@              \                 @3[Q@*Mp����?�            �i@                                  �?��]�'�?            �h@                                   @�����?             E@                                  �?��p\�?            �D@                                   �?�FVQ&�?            �@@               	                   �H@      �?              @       ������������������������       �                     @        
                        83F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?`2U0*��?             9@                                  P,@�C��2(�?             &@       ������������������������       �                      @                                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@                                83�0@      �?              @                                  �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               +                     @ގ$@�h�?a            �c@               *                    �?$G$n��?,            �R@              )                  �v7@�<ݚ�?            �F@                                `f&'@��}*_��?             ;@                                  �J@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        !       "                   �;@�z�G��?             4@        ������������������������       �                     @        #       $                   �B@��S�ۿ?
             .@       ������������������������       �                     &@        %       (                   �*@      �?             @        &       '                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �                     =@        ,       Y                 �̼6@�!>�R�?5            �T@       -       P                 �|Y=@      �?%             O@       .       ?                   �3@�zv�X�?             F@        /       >                   �2@j���� �?             1@       0       5                    '@��S���?             .@        1       2                 @3�2@z�G�z�?             @       ������������������������       �                     @        3       4                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        6       =                    �?���Q��?             $@       7       8                 P��@      �?              @        ������������������������       �                     �?        9       :                 ��!@؇���X�?             @        ������������������������       �                     @        ;       <                 `F�+@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        @       O                    �?������?             ;@       A       N                    �?�θ�?             :@       B       I                   �9@����X�?             5@       C       D                 ���@     ��?
             0@        ������������������������       �                      @        E       H                 pff@@4և���?             ,@        F       G                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        J       K                 �?�@���Q��?             @        ������������������������       �                     �?        L       M                 pf(@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        Q       X                    �?�<ݚ�?	             2@       R       W                 03�1@������?             .@       S       V                   &@�8��8��?             (@        T       U                    A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     @        Z       [                    @���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     @        ^       _                  "�b@0�z��?�?!             O@       ������������������������       �                     E@        `       a                    �?P���Q�?             4@       ������������������������       �                     &@        b       c                    $@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        e       �                 ��D:@���_�k�?           �{@       f       s                     @�T_�/��?�            `t@        g       h                    #@xdQ�m��?2            @T@        ������������������������       �                     @        i       j                 `f�)@�e���@�?.            @S@        ������������������������       �                     ?@        k       l                     �?��<b�ƥ?             G@        ������������������������       �                     �?        m       r                   �*@����?�?            �F@        n       o                    @@���N8�?             5@        ������������������������       �                     (@        p       q                   @B@�����H�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     8@        t       u                    $@�Zp���?�            �n@        ������������������������       �                     @        v       �                    �?pTjD��?�             n@        w       �                    �?b�h�d.�?1            �Q@       x       �                    �?��ɉ�?-            @P@       y       z                 ���@(N:!���?            �A@        ������������������������       �                      @        {       ~                   �5@PN��T'�?             ;@        |       }                 �y.@      �?             @       ������������������������       �                      @        ������������������������       �                      @               �                 �� @���}<S�?             7@       �       �                 �|�=@�r����?
             .@       �       �                   @@"pc�
�?             &@       �       �                 �|=@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        �       �                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y=@r�q��?             >@        �       �                  ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `3@؇���X�?             <@       �       �                 X�I@`2U0*��?             9@       �       �                 ���@ �q�q�?             8@        ������������������������       �                      @        �       �                   @'@      �?             0@       ������������������������       ��C��2(�?	             &@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@�����?j            `e@       �       �                    �?��<b�ƥ?9             W@       �       �                   �8@p�C��?8            �V@        �       �                 ���@�IєX�?             A@        �       �                 ���@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     7@        ������������������������       �        #            �L@        ������������������������       �                     �?        �       �                 `f�'@p#�����?1            �S@       �       �                 ���"@L=�m��?&            �N@       �       �                   �3@PN��T'�?              K@        �       �                 0S5 @����X�?             ,@        �       �                   �2@      �?              @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                 �|Y>@ףp=
�?             D@       �       �                 pf� @ ��WV�?             :@       ������������������������       �                     5@        �       �                 @3�!@z�G�z�?             @       �       �                   �:@�q�q�?             @        ������������������������       �                     �?        �       �                 �|Y<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 @3�@d}h���?             ,@        �       �                   �?@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     "@        �       �                   �<@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        �       �                     �?j���� �?N            �]@       �       �                 03c@V�K/��?5            �S@       �       �                   �<@��x�5��?1            @Q@        �       �                    �?ףp=
�?             4@       �       �                    �?8�Z$���?             *@        �       �                 0�HU@      �?             @       �       �                    9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 `f�D@�����H�?             "@       ������������������������       �                     @        �       �                   �;@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?Rg��J��?%            �H@       �       �                  �>@�ݏ^���?"            �F@        �       �                    �?�����?             3@        �       �                 �|�=@���Q��?             @        ������������������������       �                      @        �       �                 `f&;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @>@����X�?
             ,@       �       �                   �?@���|���?             &@        ������������������������       �                      @        �       �                   @L@�<ݚ�?             "@       �       �                 03k:@؇���X�?             @        ������������������������       �                     �?        �       �                   �C@r�q��?             @        ������������������������       �                     �?        �       �                   @G@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                    R@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�n_Y�K�?             :@        �       �                  �>@և���X�?             @        ������������������������       �                     �?        �       �                   �H@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y>@�����?             3@        ������������������������       �                     @        �       �                  x#J@և���X�?
             ,@        ������������������������       �                     @        �       �                    F@�q�q�?             "@        ������������������������       �                     @        �       �                    H@      �?             @        ������������������������       �                      @        �       �                 ���W@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @B@ףp=
�?             $@        �       �                 X�,@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �                           @z�G�z�?             D@        �       �                    �?������?
             1@        ������������������������       �                      @                                  �?X�<ݚ�?             "@                                 0@      �?             @        ������������������������       �                      @        ������������������������       �                      @                              pV�C@���Q��?             @                                �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        	                      �|�>@�LQ�1	�?             7@       
                         �?ףp=
�?             4@                                5@��S�ۿ?             .@       ������������������������       �                     "@                                 ;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                 @z�G�z�?             @                                  @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?SKE,�?WwZ�iu�?�������?�?��Aˎ��?,2_�8��?�a�a�?=��<���?��+Q��?�]�ڕ��?|���?>����?      �?      �?              �?      �?      �?      �?                      �?{�G�z�?���Q��?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?      �?        ~��	���?A����?���L�?к����?�q�q�?9��8���?B{	�%��?_B{	�%�?�$I�$I�?۶m۶m�?              �?      �?        333333�?ffffff�?      �?        �?�������?              �?      �?      �?      �?      �?      �?                      �?              �?              �?              �?+Jx���?��k���?      �?      �?��.���?�袋.��?ZZZZZZ�?�������?�������?�?�������?�������?              �?      �?      �?      �?                      �?333333�?�������?      �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?                      �?              �?B{	�%��?{	�%���?ى�؉��?�؉�؉�?�m۶m��?�$I�$I�?      �?      �?              �?n۶m۶�?�$I�$I�?      �?      �?              �?      �?              �?        �������?333333�?      �?              �?      �?              �?      �?              �?                      �?�q�q�?9��8���?�?wwwwww�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?                      �?��y��y�?�a�a�?              �?      �?              �?        �B!��?|���{�?              �?�������?ffffff�?              �?�q�q�?�q�q�?      �?                      �?�����?~������?�A2����?K�m�
��?�5?,R�?X�<ݚ�?              �?qV~B���?�cj`?      �?        ��7��M�?d!Y�B�?      �?        ��I��I�?l�l��?��y��y�?�a�a�?      �?        �q�q�?�q�q�?      �?      �?      �?              �?        Az�U6�?�-�RM�?              �?5�5��?W�W��?;��:���?_�_��?�����?�����?|�W|�W�?�A�A�?      �?        &���^B�?h/�����?      �?      �?              �?      �?        ӛ���7�?d!Y�B�?�������?�?/�袋.�?F]t�E�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?              �?      �?              �?              �?        �������?UUUUUU�?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?���Q��?{�G�z�?�������?UUUUUU�?      �?              �?      �?]t�E�?F]t�E�?      �?              �?                      �?�������?333333�?              �?      �?        �Md7��?d7��Dv�?��7��M�?d!Y�B�?��K��K�?h�h��?�?�?/�袋.�?F]t�E�?      �?                      �?      �?              �?              �?        7a~W��?�#{���?���:�?�����?&���^B�?h/�����?�m۶m��?�$I�$I�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?O��N���?;�;��?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        I�$I�$�?۶m۶m�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?        �������?ZZZZZZ�?�Z܄��?�ґ=�?�Q�g���?0�̵�?�������?�������?;�;��?;�;��?      �?      �?      �?      �?      �?                      �?              �?�q�q�?�q�q�?              �?      �?      �?              �?      �?                      �??4և���?��S�r
�?��I��I�?�[�[�?^Cy�5�?Q^Cy��?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?�m۶m��?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?              �?�������?�������?      �?      �?              �?      �?      �?      �?                      �?              �?;�;��?ى�؉��?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        Q^Cy��?^Cy�5�?      �?        �$I�$I�?۶m۶m�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?                      �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ffffff�?ffffff�?xxxxxx�?�?      �?        r�q��?�q�q�?      �?      �?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ��Moz��?Y�B��?�������?�������?�������?�?      �?        �������?UUUUUU�?              �?      �?        �������?�������?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ4�phG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM9hjh))��}�(h,h/h0M9��h2h3h4hph<�h=Kub������       �                    �?�C�"���?�           8�@              ;                     �?�#}7��?C           ��@               *                  x#J@     ��?O             `@              	                    �?z�7�Z�?,            @R@                                   �?�8��8��?             (@                                ��A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        
                          �<@�jTM��?%            �N@                                   �?      �?              @        ������������������������       �                      @                                ��iB@      �?             @        ������������������������       �                     @        ������������������������       �                     @                                   �?r�����?"            �J@                                �|�=@r�q��?             (@                                ��2>@����X�?             @                               �ܵ<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               )                  i?@� ��1�?            �D@              (                   @>@�LQ�1	�?             7@                                  A@      �?             4@                                �|Y=@�����H�?             "@        ������������������������       �                      @                                `fF<@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                !                 ��$:@���|���?
             &@        ������������������������       �                     @        "       #                 03k:@      �?              @        ������������������������       �                      @        $       '                 `f�;@�q�q�?             @       %       &                    J@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             2@        +       8                  �k@"pc�
�?#            �K@       ,       -                    �?��E�B��?            �G@       ������������������������       �                     ;@        .       /                    6@�z�G��?             4@        ������������������������       �                      @        0       1                    �?�<ݚ�?             2@        ������������������������       �                     @        2       3                 03�M@�q�q�?             (@        ������������������������       �                     @        4       5                    �?�q�q�?             @        ������������������������       �                     �?        6       7                 ��#[@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        9       :                 X�,@@      �?              @        ������������������������       �                     @        ������������������������       �                     @        <       ?                   �,@�t.��?�            �y@        =       >                    �?�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        @       �                 ���$@��ϫ��?�            �x@       A       n                 �̌@�i� ���?�            @m@        B       U                    �?P����?F            �\@        C       T                    @�J�4�?             9@       D       O                 ��@���y4F�?             3@       E       N                 X��B@      �?
             0@       F       G                    �?��S�ۿ?	             .@       ������������������������       �                     $@        H       I                 ���@z�G�z�?             @        ������������������������       �                     �?        J       M                 pff@      �?             @       K       L                 �|Y:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        P       Q                    4@�q�q�?             @        ������������������������       �                     �?        R       S                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        V       W                     @��f��?3            @V@        ������������������������       �                     @        X       ]                   @4@�~6�]�?0            @U@        Y       \                 �&�@�eP*L��?             &@       Z       [                    �?      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ^       e                    �?�MI8d�?+            �R@        _       b                 ���@H�V�e��?             A@       `       a                   �7@؇���X�?             5@        ������������������������       �                     @        ������������������������       �        
             2@        c       d                 �|Y=@�	j*D�?             *@        ������������������������       �                      @        ������������������������       �"pc�
�?             &@        f       g                 �|Y=@      �?             D@        ������������������������       �                     *@        h       m                 �&B@�+$�jP�?             ;@       i       j                 ��@�8��8��?             8@       ������������������������       �                     0@        k       l                 �|Y>@      �?              @        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        o       �                 ��) @��S�ۿ?G             ^@       p       y                 @3�@��+��<�?.            �U@       q       x                 �?�@��<b�ƥ?             G@       r       w                 �|Y=@P�Lt�<�?             C@        s       t                    �?��S�ۿ?
             .@        ������������������������       �                      @        u       v                    �?$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     7@        ������������������������       �                      @        z       {                    �?P���Q�?             D@        ������������������������       �                     @        |       �                   �3@@-�_ .�?            �B@        }       ~                    1@�q�q�?             @        ������������������������       �                     �?               �                   �2@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     ?@        �       �                    �?��hJ,�?             A@        ������������������������       �                     @        �       �                    �?�חF�P�?             ?@        ������������������������       �                     @        �       �                 ��i @���B���?             :@        ������������������������       �                     �?        �       �                 @�!@�J�4�?             9@        �       �                 pf!@      �?             (@        ������������������������       �                      @        �       �                 �|Y<@�z�G��?             $@        �       �                    6@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�=@$�q-�?             *@       ������������������������       �        
             (@        ������������������������       �                     �?        �       �                 `f�)@���|���?b            �d@        �       �                   �>@��
P��?            �A@       �       �                   �9@����X�?             5@       �       �                   �'@X�<ݚ�?             "@       �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                    4@r�q��?             @        �       �                    &@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �<@�8��8��?             (@        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �@@d}h���?	             ,@        ������������������������       �                     @        �       �                   @I@և���X�?             @        �       �                   @A@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �̌.@@i��M��?N            @`@        �       �                    �?�iʫ{�?            �J@        �       �                    �?���|���?             &@        �       �                   �2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    :@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �D@���N8�?             E@       �       �                 �|Y<@��?^�k�?            �A@        ������������������������       �                     1@        �       �                    �?�X�<ݺ?             2@        ������������������������       �                     @        �       �                     @@4և���?	             ,@       �       �                 �|�=@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �       �                   �*@؇���X�?             @       �       �                    G@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �2@և���X�?/            @S@        ������������������������       �                      @        �       �                   �E@
;&����?+            @Q@       �       �                   �C@     ��?'             P@       �       �                 �|�=@�������?%             N@       �       �                  �v6@�K��&�?            �E@       �       �                     @�û��|�?             7@        ������������������������       �                     �?        �       �                    �?8�A�0��?             6@        �       �                 ���/@�����H�?             "@        ������������������������       �                     @        �       �                 �|�;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?$�q-�?             *@        �       �                 м;4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?z�G�z�?             4@        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �;@r�q��?
             2@        �       �                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        �       �                 03�1@������?             1@        �       �                 pff/@���Q��?             @        ������������������������       �                     �?        �       �                   �0@      �?             @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�8��8��?             (@        �       �                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     @        �                           @{�����?j            �e@        �       �                    �?rEC��a�?-            �S@        �       �                     �?     ��?	             0@       �       �                    �?�eP*L��?             &@       �       �                 ��UO@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    ,@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��d��?$            �O@       ������������������������       �                     F@                                  :@�\��N��?             3@                                 *@      �?              @        ������������������������       �                     �?        ������������������������       �                     @                                 0@"pc�
�?	             &@        ������������������������       �                      @        ������������������������       �                     "@              &                   �?      �?=             X@                                �?�`���?#            �H@        	                         �?8�Z$���?	             *@       
                      83�0@����X�?             @                                &@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                 @b�2�tk�?             B@                                 �?�q�q�?	             (@                                 @z�G�z�?             @        ������������������������       �                     @                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?և���X�?             @        ������������������������       �                      @                              pf�0@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?              !                   �?      �?             8@                                 �;@X�<ݚ�?             "@                              pf�0@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        "      %                `f2@��S�ۿ?             .@        #      $                `ff/@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        '      ,                �̼6@��|�5��?            �G@        (      )                  �5@�<ݚ�?             "@        ������������������������       �                     @        *      +                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        -      6                   �?�KM�]�?             C@       .      /                   �? 7���B�?             ;@        ������������������������       �                      @        0      1                X��@@`2U0*��?             9@       ������������������������       �        	             4@        2      5                   @z�G�z�?             @       3      4                  �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        7      8                   @���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0M9KK��h2h3h4hVh<�h=Kub�������������[�e�?���I54�?~5&��?���[��?     ��?     ��?�I�&M��?�lٲe��?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�y��!�?.�u�y�?      �?      �?              �?      �?      �?              �?      �?        Dj��V��?�V�9�&�?�������?UUUUUU�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ������?������?Nozӛ��?d!Y�B�?      �?      �?�q�q�?�q�q�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?]t�E]�?F]t�E�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?              �?                      �?      �?        F]t�E�?/�袋.�?AL� &W�?�l�w6��?              �?333333�?ffffff�?      �?        �q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?                      �?      �?      �?      �?                      �?######�?�������?UUUUUU�?UUUUUU�?              �?      �?        �v��%k�?�mJ�)�?*��)���?Z��Y���?�P^Cy�?Q^Cy��?{�G�z�?�z�G��?(������?6��P^C�?      �?      �?�?�������?              �?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?���0��?��g<��?      �?        999999�?�?]t�E�?t�E]t�?      �?      �?              �?      �?              �?        ��L���?L�Ϻ��?iiiiii�?ZZZZZZ�?۶m۶m�?�$I�$I�?              �?      �?        vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?      �?      �?      �?        /�����?B{	�%��?UUUUUU�?UUUUUU�?      �?              �?      �?333333�?�������?      �?                      �?�������?�?�#�;��?w�qGܡ?��7��M�?d!Y�B�?���k(�?(�����?�������?�?      �?        �؉�؉�?;�;��?              �?      �?              �?              �?        ffffff�?�������?      �?        S�n0E�?к����?UUUUUU�?UUUUUU�?      �?        333333�?�������?              �?      �?      �?      �?        KKKKKK�?�������?      �?        �Zk����?��RJ)��?      �?        ��؉���?ى�؉��?              �?�z�G��?{�G�z�?      �?      �?      �?        ffffff�?333333�?      �?      �?      �?                      �?      �?        �؉�؉�?;�;��?      �?                      �?]t�E]�?F]t�E�?_�_��?PuPu�?�$I�$I�?�m۶m��?r�q��?�q�q�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?              �?      �?        I�$I�$�?۶m۶m�?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?              �?      �?              �?        �Z��Z��?�J��J��?
�[���?�琚`��?F]t�E�?]t�E]�?      �?      �?      �?                      �?�$I�$I�?�m۶m��?      �?                      �?��y��y�?�a�a�?_�_��?�A�A�?      �?        ��8��8�?�q�q�?      �?        n۶m۶�?�$I�$I�?]t�E�?F]t�E�?              �?      �?              �?        ۶m۶m�?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?        �$I�$I�?۶m۶m�?      �?        Y�B��?�Mozӛ�?      �?     ��?�������?�������?���)k��?��)kʚ�?8��Moz�?��,d!�?      �?        颋.���?/�袋.�?�q�q�?�q�q�?              �?      �?      �?      �?                      �?�؉�؉�?;�;��?      �?      �?              �?      �?              �?        �������?�������?      �?      �?              �?      �?        UUUUUU�?�������?۶m۶m�?�$I�$I�?              �?      �?                      �?xxxxxx�?�?�������?333333�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?      �?        v��4��?E'���?�=Q���?�0���M�?      �?      �?]t�E�?t�E]t�?�q�q�?r�q��?      �?                      �?      �?      �?              �?      �?        �������?�������?              �?      �?        EQEQ�?��뺮��?              �?y�5���?�5��P�?      �?      �?      �?                      �?/�袋.�?F]t�E�?              �?      �?              �?      �?և���X�?����S�?;�;��?;�;��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�8��8��?9��8���?UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?              �?      �?�q�q�?r�q��?UUUUUU�?�������?              �?      �?              �?        �������?�?      �?      �?      �?                      �?      �?        br1���?x6�;��?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?      �?        �k(���?(�����?	�%����?h/�����?      �?        ���Q��?{�G�z�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        F]t�E�?t�E]t�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJLxhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       h                     @��l�Qf�?�           8�@                                  �1@<W#.m��?�            �s@                                   �?���}<S�?             7@                                   3@      �?             @        ������������������������       �                      @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        	                            �?�}�+r��?             3@        
                           !@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@               %                    �?�6����?�            @r@                                   @L@PF��t<�?P            �_@                                  �? �^�@̩?K             ]@        ������������������������       �                    �E@                                    �?���(-�?1            @R@        ������������������������       �                     ?@                                  �*@@4և���?             E@                                  �'@؇���X�?	             ,@        ������������������������       �                     @                                   :@      �?              @        ������������������������       �                      @        ������������������������       �                     @                                   �?h�����?             <@                                  �E@$�q-�?	             *@       ������������������������       �                      @                                   5@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             .@        !       "                    �?�C��2(�?             &@        ������������������������       �                     @        #       $                     �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        &       W                     �?z�G�z�?f            �d@       '       V                    �?Z��:���?;            �V@       (       9                    �?t�C�#��?4            �S@        )       8                 p"�X@8����?             7@       *       1                 ��<J@j���� �?             1@       +       0                 �|�=@�����H�?             "@        ,       -                 �ܵ<@      �?             @        ������������������������       �                      @        .       /                 03SA@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        2       3                  �}S@      �?              @        ������������������������       �                     @        4       7                    �?�q�q�?             @       5       6                   �8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        :       Q                   �G@��>4և�?#             L@       ;       P                   �E@��V#�?            �E@       <       =                 ��I*@l��[B��?             =@        ������������������������       �                     @        >       E                 �|Y=@�û��|�?             7@        ?       D                   �<@����X�?             @       @       A                   �7@      �?             @        ������������������������       �                     �?        B       C                 `f�D@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        F       O                   �B@      �?             0@       G       N                    B@���|���?             &@       H       M                   �D@�z�G��?             $@       I       L                 `fF<@      �?              @       J       K                 X�,@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        R       S                   �J@�n_Y�K�?
             *@        ������������������������       �                     @        T       U                    R@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        X       g                   �*@@-�_ .�?+            �R@       Y       ^                   �)@�����?             E@        Z       ]                    &@���N8�?             5@       [       \                    5@@4և���?             ,@        ������������������������       �z�G�z�?             @        ������������������������       �                     "@        ������������������������       �                     @        _       `                 �|�<@؇���X�?             5@        ������������������������       �                     $@        a       b                 �|�=@���!pc�?             &@        ������������������������       �                     �?        c       f                   �A@z�G�z�?             $@       d       e                    @@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @@        i       
                  �C@      �?�            �x@       j       �                    �?����n�?�            �v@        k       �                   �<@��k��?D            �Z@       l       �                    @     8�?&             P@       m       �                    �?�U���?%             O@       n       o                 ��@�eP*L��?            �@@        ������������������������       �                     @        p       u                    �?�q�q�?             ;@        q       r                   �,@      �?             @        ������������������������       �                      @        s       t                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        v       }                   �9@��+7��?             7@       w       x                  �#@�����H�?	             2@       ������������������������       �                     (@        y       |                    4@�q�q�?             @       z       {                 �y�+@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ~       �                 �?�@z�G�z�?             @              �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @J�8���?             =@        �       �                    �?      �?              @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �*@���N8�?             5@        ������������������������       �                     @        �       �                    5@�IєX�?             1@       ������������������������       �                     *@        �       �                    :@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?0,Tg��?             E@       �       �                 м[8@؇���X�?            �A@       �       �                    �?�C��2(�?            �@@        ������������������������       �                     �?        �       �                   �>@      �?             @@       �       �                    �?`2U0*��?             9@       ������������������������       �                     2@        �       �                 pf�$@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?؇���X�?             @       �       �                 03�1@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y=@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?    �7�?�             p@       �       �                   �B@>����?�            @k@       �       �                    �?�g��?�            �j@        �       �                   �:@��R[s�?            �A@        �       �                 ��y@���|���?             &@        ������������������������       �                      @        �       �                 �&�)@�<ݚ�?             "@       ������������������������       �                     @        �       �                 �0@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �|Y=@�8��8��?             8@        �       �                   �<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���@P���Q�?             4@        ������������������������       �                     $@        �       �                   @@ףp=
�?             $@       �       �                 �|�=@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �T)D@�����H�?w            �f@       �       �                 @3�@���i�V�?u             f@       �       �                    �?      �?B             Z@        �       �                  s�@�t����?
             1@        ������������������������       �                     @        �       �                 ��(@8�Z$���?             *@       ������������������������       �"pc�
�?             &@        ������������������������       �                      @        �       �                   �?@�=C|F�?8            �U@       �       �                   �8@�����?/            �R@        �       �                 �?�@b�h�d.�?            �A@       �       �                   �7@ܷ��?��?             =@       ������������������������       �                     6@        �       �                 `fF@և���X�?             @        �       �                 �&b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �4@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �&B@ ���J��?            �C@        �       �                 �|�;@      �?              @        ������������������������       �                     @        �       �                 �|Y>@�q�q�?             @       �       �                 pf�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ?@        �       �                 03�@�	j*D�?	             *@        ������������������������       �                     @        �       �                   �@      �?              @        ������������������������       �                     �?        �       �                 �?�@և���X�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        �       �                   �:@�X�<ݺ?3             R@        ������������������������       �                     <@        �       �                 03�6@�C��2(�?             F@       �       �                   �;@@4և���?             E@        ������������������������       �                      @        �       �                 ���"@�(\����?             D@        ������������������������       �                     5@        �       �                    �?�}�+r��?             3@        ������������������������       �                     @        �       �                 �|�=@      �?             0@       ������������������������       �                     (@        �       �                 ��)@      �?             @       �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�I�w�"�?             C@        �       �                 ��y&@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?     ��?             @@        ������������������������       �                     �?               	                   #@�חF�P�?             ?@                                 @�n_Y�K�?             *@                                �?      �?              @       ������������������������       �                     @                              pf�@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                              `f�9@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     A@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������}<����?�/���?��	��	�?�����?d!Y�B�?ӛ���7�?      �?      �?              �?      �?      �?              �?      �?        (�����?�5��P�?�������?�������?      �?                      �?              �?�ܹs���?�#F��?�@ �?�������?a���{�?5�rO#,�?              �?�P�B�
�?��իW��?              �?�$I�$I�?n۶m۶�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?�$I�$I�?�m۶m��?;�;��?�؉�؉�?              �?�������?�������?              �?      �?                      �?F]t�E�?]t�E�?              �?      �?      �?              �?      �?        �������?�������?�\��\��?TFeTFe�?��td�@�?��7a~�?d!Y�B�?8��Moz�?�������?ZZZZZZ�?�q�q�?�q�q�?      �?      �?      �?              �?      �?              �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        ۶m۶m�?I�$I�$�?eMYS֔�?6eMYS��?���=��?GX�i���?      �?        ��,d!�?8��Moz�?�m۶m��?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?F]t�E�?]t�E]�?333333�?ffffff�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?                      �?      �?        ى�؉��?;�;��?              �?�m۶m��?�$I�$I�?      �?                      �?      �?        S�n0E�?к����?=��<���?�a�a�?��y��y�?�a�a�?n۶m۶�?�$I�$I�?�������?�������?      �?              �?        ۶m۶m�?�$I�$I�?      �?        F]t�E�?t�E]t�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?      �?��{�?�?���	���?"5�x+��?oe�Cj��?     ��?      �?c�1��?�9�s��?t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?      �?                      �?zӛ����?Y�B��?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?333333�?�������?              �?      �?              �?        �������?�������?      �?      �?              �?      �?                      �?�rO#,��?|a���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �������?333333�?      �?                      �?�a�a�?��y��y�?              �?�?�?      �?              �?      �?              �?      �?                      �?1�0��?�y��y��?�$I�$I�?۶m۶m�?F]t�E�?]t�E�?      �?              �?      �?{�G�z�?���Q��?              �?�$I�$I�?۶m۶m�?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?             ��?     ��?ش�,�M�?�,�M���?��U��?�=��C�?X|�W|��?PuPu�?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?ffffff�?�������?      �?        �������?�������?�������?�������?      �?      �?      �?              �?        �q�q�?�q�q�?颋.���?�袋.��?      �?      �?<<<<<<�?�?      �?        ;�;��?;�;��?/�袋.�?F]t�E�?      �?        �C��:��?J��/�?�Ϻ���?v�)�Y7�?;��:���?_�_��?��=���?a���{�?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        ��-��-�?�A�A�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        vb'vb'�?;�;��?      �?              �?      �?              �?�$I�$I�?۶m۶m�?      �?              �?      �?��8��8�?�q�q�?      �?        ]t�E�?F]t�E�?n۶m۶�?�$I�$I�?              �?333333�?�������?      �?        �5��P�?(�����?      �?              �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?              �?      �?      �?                      �?              �?����k�?�5��P�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?        �Zk����?��RJ)��?;�;��?ى�؉��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW��8hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       b                    �?H���I�?�           8�@               K                   �>@���N8�?�            �o@              :                    �?���f+�?i            `e@              3                 `v�5@�xK���?R            `a@                                   @��j���?5            �T@                                   1@     ��?	             0@              
                   �9@@4և���?             ,@               	                    )@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                 ��@�d�K���?,            �P@                                   �?z�G�z�?            �A@                               �|�9@�KM�]�?             3@        ������������������������       �                      @                                ���@"pc�
�?	             &@        ������������������������       �                      @        ������������������������       �                     "@                                 s@     ��?             0@        ������������������������       �                     @                                pff@�q�q�?             (@                                �|Y:@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                ���@z�G�z�?             @        ������������������������       �                      @                                   4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               "                    @      �?             @@                !                 ��*4@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        #       ,                   �9@�+e�X�?             9@       $       +                    3@�IєX�?             1@        %       &                    �?      �?              @        ������������������������       �                     @        '       *                    �?z�G�z�?             @       (       )                 �y�+@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        -       .                    �?      �?              @        ������������������������       �                     �?        /       2                 �|Y=@����X�?             @       0       1                    <@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        4       5                    �?h�����?             L@       ������������������������       �                     C@        6       7                 03�7@�����H�?             2@        ������������������������       �                      @        8       9                 039@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ;       >                     @     ��?             @@        <       =                    @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ?       F                 �̼6@���!pc�?             6@        @       E                    @X�<ݚ�?             "@       A       D                   �/@      �?              @        B       C                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        G       H                 ��T?@$�q-�?
             *@        ������������������������       �                     @        I       J                 ��p@@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        L       ]                     @�
��P�?1            @T@       M       R                    �? >�֕�?*            �Q@        N       Q                    �?�8��8��?	             (@       O       P                 8��J@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        S       V                   �'@�8���?!             M@        T       U                   �J@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        W       X                     �?`Ql�R�?            �G@        ������������������������       �                     2@        Y       Z                   �B@XB���?             =@       ������������������������       �        	             2@        [       \                   �C@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ^       _                    �?���|���?             &@        ������������������������       �                     @        `       a                   �B@      �?              @        ������������������������       �                     @        ������������������������       �                     @        c       �                 03s/@��`��?           �|@       d       s                    �?�hrF��?�            ps@        e       j                   �6@>A�F<�?             C@        f       i                 ��}@z�G�z�?             @       g       h                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        k       l                     @�C��2(�?            �@@        ������������������������       �                      @        m       n                 ���@��a�n`�?             ?@        ������������������������       �                     ,@        o       r                 �|�=@@�0�!��?	             1@       p       q                   @@���!pc�?             &@       ������������������������       �և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        t       �                     @�o�ا?�?�            q@        u       v                 ��"@6uH���?!             O@        ������������������������       �                      @        w       x                     �?P���Q�?              N@        ������������������������       �                     $@        y       �                    �? "��u�?             I@       z                           4@=QcG��?            �G@        {       |                   �2@�q�q�?             @        ������������������������       �                     �?        }       ~                   �'@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                   �C@��Y��]�?            �D@       ������������������������       �                     >@        �       �                   @F@�C��2(�?             &@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �?�@P�S�L�?�            `j@       �       �                   �<@�-.�1a�?F            �^@        ������������������������       �                     K@        �       �                    �?��.N"Ҭ?(            @Q@        �       �                  s�@�KM�]�?             3@        ������������������������       �                     @        �       �                 ��(@؇���X�?             ,@       �       �                 �|Y=@8�Z$���?
             *@        ������������������������       �                     �?        �       �                 X��A@�8��8��?	             (@       ������������������������       �ףp=
�?             $@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     I@        �       �                 @3�@h�V���?<             V@        �       �                   �?@      �?             (@        �       �                    :@���Q��?             @       �       �                   �4@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �A@؇���X�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                    &@�˹�m��?4             S@        ������������������������       �                     �?        �       �                    �?��S�ۿ?3            �R@        ������������������������       �                     @        �       �                    �?D��*�4�?/            @Q@       �       �                 ��) @�U�=���?-            �P@        �       �                    3@�g�y��?             ?@        ������������������������       �      �?              @        ������������������������       �                     =@        �       �                   �<@(N:!���?            �A@        ������������������������       �                     .@        �       �                 �|Y=@z�G�z�?             4@        ������������������������       �                     �?        �       �                    ?@�S����?             3@        �       �                 �|�=@      �?             (@       �       �                 pf� @"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @      �?a            �b@        �       �                     @���Q��?
             .@        ������������������������       �                     @        �       �                 @3�4@�eP*L��?             &@        ������������������������       �                     @        �       �                 ��A>@؇���X�?             @        ������������������������       �                     @        �       �                 ���A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �                         @I@���y4F�?W            �`@       �                         �G@�G�.o�?J            @[@       �       �                     �?���q��?F            �Y@        �       �                    �?����X�?#             L@        �       �                    �?�ՙ/�?             5@       �       �                  �>@      �?             0@       �       �                    B@�q�q�?             "@       �       �                 ��";@և���X�?             @        ������������������������       �                     �?        �       �                 �|�=@�q�q�?             @       �       �                 �ܵ<@      �?             @        ������������������������       �                     �?        �       �                 ��2>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �4@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @       �       �                 0�HU@      �?             @       �       �                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?4�2%ޑ�?            �A@        ������������������������       �                      @        �       �                    D@r٣����?            �@@       �       �                   �;@D�n�3�?             3@        ������������������������       �                      @        �       �                 �|Y>@ҳ�wY;�?             1@       �       �                 �|Y=@�θ�?	             *@        �       �                   �<@z�G�z�?             @       �       �                 ��iB@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   `@@      �?              @        �       �                 `fF<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    B@      �?             @        ������������������������       �                      @        �       �                 03�Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                 �T�I@��E�B��?#            �G@       �       �                   �7@�˹�m��?             C@        �       �                    6@r�q��?             2@       �       �                    $@�t����?             1@        ������������������������       �                     �?        �       �                    �?      �?
             0@       �       �                    �?�����H�?             "@        �       �                   �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �                          �?�q�q�?             "@       �       �                     @      �?             @        ������������������������       �                      @                                  ;@      �?             @        ������������������������       �                      @                                 >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     8@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������Q�Ȟ���?^-n����?��y��y�?�a�a�?m%���V�?Im%����?4,�T�w�?���j��?o4u~�!�?�e�@	o�?      �?      �?�$I�$I�?n۶m۶�?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?        ����?�rv��?�������?�������?(�����?�k(���?              �?F]t�E�?/�袋.�?      �?                      �?      �?      �?              �?�������?�������?�$I�$I�?۶m۶m�?              �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�$I�$I�?۶m۶m�?              �?      �?        R���Q�?���Q��?�?�?      �?      �?      �?        �������?�������?      �?      �?              �?      �?              �?              �?              �?      �?      �?        �$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?�$I�$I�?�m۶m��?              �?�q�q�?�q�q�?              �?�������?�������?      �?                      �?      �?      �?�������?�������?      �?                      �?F]t�E�?t�E]t�?�q�q�?r�q��?      �?      �?�������?�������?      �?                      �?              �?              �?�؉�؉�?;�;��?      �?        �������?UUUUUU�?              �?      �?        ��ӭ�a�?������?�A�A�?��+��+�?UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?                      �?              �?a���{�?j��FX�?F]t�E�?/�袋.�?              �?      �?        W�+�ɕ?}g���Q�?              �?�{a���?GX�i���?              �?F]t�E�?]t�E�?      �?                      �?]t�E]�?F]t�E�?      �?              �?      �?              �?      �?        |&�{&��?f�f��?��U()��?e#S���?������?Cy�5��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?]t�E�?F]t�E�?      �?        �s�9��?�c�1Ƹ?      �?        ZZZZZZ�?�������?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?              �?        �����?���?k���Zk�?��RJ)��?              �?ffffff�?�������?      �?        �G�z�?���Q��?x6�;��?AL� &W�?UUUUUU�?UUUUUU�?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?        8��18�?������?      �?        ]t�E�?F]t�E�?      �?      �?      �?              �?        `�
��T�?JQ/#��?{����z�?�h
���?      �?        �3J���?ہ�v`��?�k(���?(�����?      �?        ۶m۶m�?�$I�$I�?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?�������?�������?      �?              �?              �?        �袋.��?/�袋.�?      �?      �?333333�?�������?      �?      �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?��P^Cy�?^Cy�5�?              �?�������?�?      �?        ہ�v`��?)�3J���?�M6�d��?e�M6�d�?��{���?�B!��?      �?      �?      �?        |�W|�W�?�A�A�?      �?        �������?�������?              �?(������?^Cy�5�?      �?      �?/�袋.�?F]t�E�?              �?      �?                      �?      �?              �?              �?      �?�������?333333�?              �?t�E]t�?]t�E�?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        6��P^C�?(������?z|���?��p�?�e�@*�?ch���V�?�m۶m��?�$I�$I�?�<��<��?�a�a�?      �?      �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?      �?      �?      �?      �?                      �?              �?              �?      �?        �������?�A�A�?      �?        >���>�?|���?l(�����?(������?              �?�������?�������?ى�؉��?�؉�؉�?�������?�������?      �?      �?              �?      �?              �?              �?      �?      �?      �?      �?                      �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        �l�w6��?AL� &W�?��P^Cy�?^Cy�5�?�������?UUUUUU�?<<<<<<�?�?              �?      �?      �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��UhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       ^                    �?e�L��?�           8�@               %                     @��,?S�?�            @n@                                  @@2����?Z            �a@        ������������������������       �                      @               $                 03�<@�%IM��?Y            �a@               #                    �?�חF�P�?+             O@              "                 03[;@�GN�z�?             F@                                 �2@��s����?             E@       	       
                    �?ȵHPS!�?             :@        ������������������������       �                     @                                   L@R���Q�?             4@                                 �9@�KM�]�?             3@                                  �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                `f�)@�IєX�?             1@        ������������������������       �                     @                                  �B@ףp=
�?	             $@       ������������������������       �                     @                                  �C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                    �?     ��?	             0@        ������������������������       �                      @                                   �?X�Cc�?             ,@        ������������������������       �                     �?                                  �7@�n_Y�K�?             *@                                   ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                !                    D@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �        .            �S@        &       ]                 ��Y7@�fSO��?@            �X@       '       \                    @��Q���?5             T@       (       [                   @B@$��m��?4            �S@       )       6                    �?��M��?1            �Q@        *       +                 ���@      �?             @@        ������������������������       �                     �?        ,       -                    �?��a�n`�?             ?@       ������������������������       �                     2@        .       5                 `�@1@�θ�?             *@       /       0                    &@      �?             @        ������������������������       �                     �?        1       2                 03�-@���Q��?             @        ������������������������       �                      @        3       4                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        7       Z                    @@�e����?            �C@       8       Q                   �;@��J�fj�?            �B@       9       P                   �9@d��0u��?             >@       :       M                   �6@
j*D>�?             :@       ;       L                   �5@�q�q�?             5@       <       K                    �?     ��?             0@       =       J                   �3@��S���?
             .@       >       E                    �?�n_Y�K�?             *@       ?       D                   �2@���Q��?             $@       @       A                 P��@�q�q�?             @        ������������������������       �                     �?        B       C                    '@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        F       G                    @�q�q�?             @        ������������������������       �                     �?        H       I                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        N       O                 pf�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        R       S                 �|Y=@����X�?             @        ������������������������       �                     @        T       U                 pf�'@      �?             @        ������������������������       �                     �?        V       Y                    �?�q�q�?             @       W       X                 �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@        _       �                     �?�Y����?0           P}@        `       �                   @J@���q��?D            �]@       a       �                   �G@��C����?9            �W@       b       c                 03:@�;u�,a�?2            �S@        ������������������������       �                     &@        d       �                    �?      �?+             Q@       e       ~                   �E@�ݜ����?%            �M@       f       }                 �U�X@Tt�ó��?            �H@       g       x                  x#J@���Q��?            �F@       h       w                   �@@�g�y��?             ?@       i       p                    �?����X�?             5@        j       o                   @@@�q�q�?             (@       k       l                   �<@r�q��?             @        ������������������������       �                     @        m       n                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        q       v                 `fF<@�����H�?             "@        r       s                 03k:@      �?             @        ������������������������       �                     �?        t       u                 �|�<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        y       z                    �?؇���X�?             ,@        ������������������������       �                      @        {       |                    7@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @               �                    �?ףp=
�?             $@        ������������������������       �                      @        �       �                  I>@      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                    9@�q�q�?             "@        ������������������������       �                     @        �       �                 @��v@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                 xCQ@      �?             0@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   @I@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �H@ףp=
�?             $@        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �? �q�q�?             8@       �       �                 ���=@P���Q�?	             4@        ������������������������       �                     &@        �       �                   �R@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���@�,u�3�?�            �u@        ������������������������       �                    �@@        �       �                 ��@\_�}d�?�            �s@        ������������������������       �                     �?        �       �                    �?���!���?�            �s@       �       �                 �?$@���P��?�            0q@        �       �                  ��@���-T��?,             O@       �       �                    �? >�֕�?            �A@        �       �                   �6@�r����?             .@        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �                     4@        �       �                    8@������?             ;@        ������������������������       �                     @        �       �                    �?�q�q�?             5@       �       �                 �|Y=@����X�?             ,@        ������������������������       �                      @        �       �                 X��A@r�q��?
             (@       ������������������������       ��<ݚ�?             "@        ������������������������       �                     @        �       �                 �|Y?@և���X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        �       �                    �?4Č���?�            �j@        �       �                     @���N8�?             5@        ������������������������       �                      @        �       �                    �?�n_Y�K�?             *@       �       �                 �� @      �?              @        ������������������������       �                     @        �       �                   �:@z�G�z�?             @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `3@z�G�z�?             @       ������������������������       �                     @        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �3@      �?|             h@        �       �                   �1@r�q��?             8@        ������������������������       �                     "@        �       �                     @������?             .@        �       �                    &@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @���N8�?k             e@        �       �                   �*@��(\���?             D@       �       �                 �|Y=@�����H�?             ;@        ������������������������       �        	             (@        �       �                 �|Y>@z�G�z�?
             .@        ������������������������       �                     �?        �       �                   �C@؇���X�?	             ,@        ������������������������       �                     @        �       �                 `f�)@�<ݚ�?             "@        ������������������������       �                     �?        �       �                    G@      �?              @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �        
             *@        �       �                 �?�@     8�?N             `@        ������������������������       �                     G@        �       �                 @3�@0��P�?7            �T@        �       �                   �?@�<ݚ�?             "@       �       �                   �=@�q�q�?             @       �       �                   �4@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �;@���(-�?/            @R@        �       �                   �:@ףp=
�?             4@       �       �                    9@�}�+r��?             3@       ������������������������       �        	             .@        �       �                 �!J@@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�=@�O4R���?"            �J@       ������������������������       �                     A@        �       �                    ?@�}�+r��?             3@        �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        �                            @���?            �D@        �       �                   �:@���|���?             &@        �       �                   `6@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 pV�C@؇���X�?             @       �       �                    �?      �?             @       �       �                    0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 @z�G�z�?             >@             	                   0@d}h���?             <@                                 �?      �?              @                              ��y&@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 +@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        
                         �?ףp=
�?             4@        ������������������������       �                     (@                              �̌4@      �?              @        ������������������������       �                     �?                              ��T?@؇���X�?             @        ������������������������       �                     @                                 @      �?             @                                  @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������v�S(��?��X��?����|��?�ˠT�?-)D�{�?�7�P�?      �?        I8�y�'�?�X����?��RJ)��?�Zk����?]t�E�?�袋.��?�a�a�?z��y���?�؉�؉�?��N��N�?              �?333333�?333333�?(�����?�k(���?      �?      �?              �?      �?        �?�?              �?�������?�������?              �?      �?      �?      �?                      �?      �?              �?      �?              �?�m۶m��?%I�$I��?              �?ى�؉��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?333333�?ffffff�?              �?      �?              �?                      �?              �?�v�ļ�?w�ļ�!�?�������?333333�?vb'vb'�?�N��N��?�@�6�?��.�d��?      �?      �?      �?        �c�1Ƹ?�s�9��?              �?�؉�؉�?ى�؉��?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�A�A�?�-��-��?к����?�"�u�)�?wwwwww�?DDDDDD�?;�;��?b'vb'v�?UUUUUU�?UUUUUU�?      �?      �?�������?�?ى�؉��?;�;��?�������?333333�?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?              �?�������?�������?              �?      �?                      �?�m۶m��?�$I�$I�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?      �?                      �?      �?        ��¯�D�?���@���?�\�\�?��F��F�?#�X��?��%N��?ud�@T:�?7a~W��?      �?              �?      �?�}ylE��?W'u_�?/�����?h�����?�������?333333�?�B!��?��{���?�$I�$I�?�m۶m��?�������?�������?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?�q�q�?�q�q�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?�������?      �?                      �?      �?        �������?�������?      �?              �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?      �?      �?      �?        �������?333333�?      �?                      �?�������?�������?              �?      �?      �?      �?                      �?�������?UUUUUU�?ffffff�?�������?      �?        �q�q�?�q�q�?      �?                      �?      �?        yc���?5��g�?      �?        �y��C�?t0�O�?              �?��	�Z�?T:�g *�?����{��?4B�!4�?[k���Z�?�RJ)���?��+��+�?�A�A�?�������?�?              �?      �?              �?        B{	�%��?{	�%���?      �?        UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?9��8���?�q�q�?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?        �Xޫ-r�?}8��n�?�a�a�?��y��y�?      �?        ;�;��?ى�؉��?      �?      �?              �?�������?�������?      �?      �?      �?                      �?      �?        �������?�������?      �?              �?      �?              �?      �?              �?      �?�������?UUUUUU�?      �?        wwwwww�?�?�$I�$I�?۶m۶m�?              �?      �?              �?      �?              �?      �?        ��y��y�?�a�a�?�������?333333�?�q�q�?�q�q�?      �?        �������?�������?              �?۶m۶m�?�$I�$I�?      �?        9��8���?�q�q�?      �?              �?      �?      �?      �?      �?              �?             ��?      �?      �?        ���|�?8��18�?9��8���?�q�q�?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��իW��?�P�B�
�?�������?�������?�5��P�?(�����?      �?              �?      �?      �?                      �?              �?:�&oe�?�x+�R�?      �?        �5��P�?(�����?      �?      �?      �?                      �?      �?        28��1�?8��18�?]t�E]�?F]t�E�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?      �?              �?      �?              �?              �?        �������?�������?I�$I�$�?۶m۶m�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?              �?      �?        �������?�������?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��DphG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       j                     @@t]q�V�?�           8�@                                   �?�So���?�            �s@                                   6@���}��?S            �`@                                  @4@4?,R��?             B@                               ���*@l��\��?             A@                                 �B@      �?             8@       ������������������������       �        	             1@               	                    D@և���X�?             @        ������������������������       �                      @        
                          �J@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @                                   @��4+̰�?>            @X@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �H@ r���?<            �W@       ������������������������       �        4             T@                                �DD@�r����?             .@                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@               1                    �?�������?u            �f@               .                     �?      �?             D@              +                    �?���@M^�?             ?@              &                 X�,@@�G��l��?             5@              %                  �}S@���!pc�?             &@                                �ܵ<@և���X�?             @        ������������������������       �                      @        !       "                  Y>@���Q��?             @        ������������������������       �                      @        #       $                 �|Y<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        '       *                 @�pX@z�G�z�?             $@       (       )                   @J@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ,       -                   �7@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        /       0                    (@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        2       Q                 `ff:@������?\            �a@       3       4                     �?$�q-�?6            �S@        ������������������������       �                     @        5       J                   �7@@�j;��?0            �Q@       6       7                    @0G���ջ?%             J@        ������������������������       �                     @        8       I                   �F@=QcG��?!            �G@       9       H                    �?�˹�m��?             C@       :       =                    &@�8��8��?             B@        ;       <                   �5@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        >       G                   @D@ 	��p�?             =@       ?       @                 `fF)@ 7���B�?             ;@        ������������������������       �                      @        A       F                    1@�}�+r��?             3@       B       C                 �|Y<@�X�<ݺ?             2@       ������������������������       �                     $@        D       E                 �|�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     "@        K       P                    :@�S����?             3@       L       M                    �?@�0�!��?
             1@       ������������������������       �                     &@        N       O                   �3@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        R       g                    �?�BE����?&             O@       S       ^                   �>@�e�,��?#            �M@        T       ]                     �?�q�q�?             8@       U       Z                   �J@���!pc�?             6@       V       W                   �C@      �?             0@       ������������������������       �                     "@        X       Y                   @G@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        [       \                 `fF<@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        _       d                 ���[@�#-���?            �A@       `       c                   �D@      �?             @@        a       b                   �B@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        e       f                 X��C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        h       i                 `�fK@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        k       �                    �?�y���?�            �x@        l       �                    �?z�):���?D             Y@       m       r                    �?����"�?'             M@        n       o                 �&�)@д>��C�?             =@       ������������������������       �                     2@        p       q                  S�-@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        s       �                 ��&@�f7�z�?             =@       t       {                   �5@�d�����?             3@        u       z                   �4@և���X�?             @       v       y                   �3@      �?             @        w       x                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        |                           ;@�8��8��?	             (@       }       ~                   �9@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�;@�z�G��?             $@        �       �                 @3�,@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @���N8�?             E@        ������������������������       �                      @        �       �                    @z�G�z�?             D@       �       �                 �|Y>@     ��?             @@       �       �                    :@��� ��?             ?@       �       �                    �?�<ݚ�?             2@        ������������������������       �                     @        �       �                    1@������?             .@       �       �                    @�C��2(�?             &@        �       �                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���9@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     �?        �       �                  18@      �?              @        ������������������������       �                      @        �       �                 ��p@@r�q��?             @        �       �                 ��A>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                  s�@��� ��?�            �r@        �       �                    �?��.N"Ҭ?'            @Q@        �       �                 ���@��S�ۿ?             >@       ������������������������       �        	             3@        �       �                    �?"pc�
�?             &@       �       �                   �5@      �?              @        ������������������������       �                     �?        �       �                 �|=@؇���X�?             @        ������������������������       �                      @        �       �                 �|�=@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        �       �                    �?6�G�1��?�            �l@        �       �                    �?z�G�z�?             @       �       �                 8#8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?>4և�z�?�             l@        �       �                 �|Y=@��S���?
             .@        �       �                 ؼC1@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|Y?@�<ݚ�?             "@       �       �                  S�'@����X�?             @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�'����?�             j@       �       �                    �?���O1��?m            �d@        �       �                 �|Y=@      �?	             (@        ������������������������       �                     �?        �       �                 X��A@"pc�
�?             &@       �       �                 `f�/@�<ݚ�?             "@       ������������������������       �����X�?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �<@��2(&�?d            @c@       �       �                 �?�@��p\�?7            �T@        ������������������������       �                     :@        �       �                   �2@ �Cc}�?#             L@        �       �                   �1@���!pc�?	             &@       �       �                 pf� @�<ݚ�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        �       �                 ��Y @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�!@��S�ۿ?            �F@        �       �                 @3�@�LQ�1	�?             7@        �       �                   �4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �:@�KM�]�?
             3@       �       �                 0S5 @�X�<ݺ?	             2@       �       �                   �4@ףp=
�?             $@        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@        �       �                 @3�@�q�q�?-             R@        �       �                 �?�@��>4և�?             <@       �       �                   �@�d�����?             3@        �       �                   @@@      �?             $@       �       �                   �?@X�<ݚ�?             "@       �       �                 �|Y>@      �?              @       ������������������������       �և���X�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �?@�q�q�?             "@        ������������������������       �                     @        �       �                   �A@      �?             @       ������������������������       �      �?             @        ������������������������       �      �?              @        �       �                 �|Y=@�C��2(�?             F@        ������������������������       �                     @        �       �                 �|�=@��Y��]�?            �D@       ������������������������       �                     9@        �       �                 ��)"@      �?             0@       ������������������������       �        	             (@        �       �                 ���'@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?Du9iH��?            �E@        ������������������������       �                      @        �                           0@��p\�?            �D@        �       �                 `ff.@�<ݚ�?             "@       �       �                    &@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                              ��T?@      �?             @@       ������������������������       �        	             1@                              ���A@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������
���?�;����?��܂`��?������?���̮?4�τ?�?r�q��?�8��8��?�������?------�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?                      �?      �?         tT����?_\����?      �?      �?              �?      �?        �X�0Ҏ�?9�{n�S�?              �?�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?      �?�s�9��?�c�1��?��y��y�?1�0��?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?�q�q�?�q�q�?              �?      �?              �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        B�A��?�������?�؉�؉�?;�;��?      �?        w�'�K�?H���@��?vb'vb'�?�؉�؉�?      �?        x6�;��?AL� &W�?��P^Cy�?^Cy�5�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        ������?�{a���?	�%����?h/�����?      �?        �5��P�?(�����?��8��8�?�q�q�?      �?              �?      �?              �?      �?              �?              �?      �?      �?              �?        (������?^Cy�5�?ZZZZZZ�?�������?      �?              �?      �?              �?      �?              �?        )��RJ)�?���Zk��?�pR���?_[4��?UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?      �?      �?              �?�$I�$I�?۶m۶m�?      �?                      �?�������?UUUUUU�?      �?                      �?      �?        �A�A�?_�_�?      �?      �?�q�q�?�q�q�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�큍��?
H�Ʌ��?H�z�G�?q=
ףp�?�i��F�?	�=����?|a���?a���{�?              �?]t�E�?t�E]t�?      �?                      �?O#,�4��?a���{�?Cy�5��?y�5���?۶m۶m�?�$I�$I�?      �?      �?      �?      �?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?                      �?      �?        333333�?ffffff�?      �?      �?              �?      �?                      �?�a�a�?��y��y�?              �?�������?�������?      �?      �?�{����?�B!��?9��8���?�q�q�?      �?        wwwwww�?�?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?              �?                      �?      �?      �?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��Ug��?7`��c.�?�3J���?ہ�v`��?�������?�?      �?        /�袋.�?F]t�E�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?      �?      �?              �?              �?        =i����?
�[|=�?�������?�������?      �?      �?              �?      �?                      �?I�$I�$�?۶m۶m�?�?�������?UUUUUU�?�������?              �?      �?        9��8���?�q�q�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        !ղ���?|�4�/��?P�M�_�?���ˊ��?      �?      �?              �?/�袋.�?F]t�E�?9��8���?�q�q�?�m۶m��?�$I�$I�?      �?              �?        ��.���?t�E]t�?�]�ڕ��?��+Q��?      �?        %I�$I��?۶m۶m�?F]t�E�?t�E]t�?9��8���?�q�q�?      �?      �?      �?              �?      �?              �?      �?        �������?�?��Moz��?Y�B��?      �?      �?              �?      �?        �k(���?(�����?��8��8�?�q�q�?�������?�������?      �?      �?      �?              �?                      �?      �?        UUUUUU�?�������?۶m۶m�?I�$I�$�?Cy�5��?y�5���?      �?      �?�q�q�?r�q��?      �?      �?۶m۶m�?�$I�$I�?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?      �?      �?]t�E�?F]t�E�?              �?8��18�?������?      �?              �?      �?      �?              �?      �?              �?      �?        qG�w��?w�qGܱ?      �?        �]�ڕ��?��+Q��?9��8���?�q�q�?      �?      �?              �?      �?                      �?      �?      �?      �?        �������?�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ%�[6hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������                           @��l�Qf�?�           8�@                                    �?��k=.��?            �G@                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @                                   @�T|n�q�?            �E@                                    @���Q��?
             .@        ������������������������       �                     @        	       
                    �?      �?              @        ������������������������       �                      @                                (C45@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                   @h�����?             <@                                ���7@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             6@               ^                    �?F�O�Ko�?�           ��@               K                   @C@^��e��?�            �j@                                   @��P���?j            �d@                                  6@��K2��?8            �W@                                   �?�X�<ݺ?             2@        ������������������������       �                     @                                  @4@$�q-�?	             *@       ������������������������       �                     &@                                   ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        +             S@               .                    �?      �?2            �Q@                '                 �&�)@����"�?             =@       !       &                    �?      �?             4@       "       #                    �?�t����?             1@        ������������������������       �                      @        $       %                 ���@�r����?             .@        ������������������������       �                      @        ������������������������       �        
             *@        ������������������������       �                     @        (       )                    5@�q�q�?             "@        ������������������������       �                     @        *       -                    �?      �?             @       +       ,                 ���0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        /       0                 pf�@v�2t5�?            �D@        ������������������������       �                     @        1       >                   �:@p�ݯ��?             C@       2       9                    �?�+e�X�?             9@       3       8                   �3@�t����?             1@        4       7                   �2@      �?             @       5       6                 �y�+@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        :       ;                    �?      �?              @        ������������������������       �                      @        <       =                 ���7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ?       J                    @�n_Y�K�?             *@       @       I                 `fV6@�q�q�?
             (@       A       D                    �?�<ݚ�?             "@       B       C                 ��1@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        E       F                    <@z�G�z�?             @        ������������������������       �                     @        G       H                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        L       ]                    @`�(c�?            �H@       M       P                    �?���y4F�?             C@        N       O                 ��A@z�G�z�?
             .@        ������������������������       �                     @        ������������������������       �        	             (@        Q       V                   @.@��<b���?             7@        R       U                    G@�q�q�?             @       S       T                   @%@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        W       X                     �?�IєX�?             1@       ������������������������       �                      @        Y       \                    G@�����H�?             "@       Z       [                   �6@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        _       �                     �?���av��?"           0|@        `       y                    �?4�E��
�?>             Z@        a       b                 `f&;@�g�y��?             ?@        ������������������������       �                      @        c       j                 �D�G@l��[B��?             =@        d       i                  Y>@���!pc�?             &@        e       f                 ���<@���Q��?             @        ������������������������       �                     �?        g       h                 X��E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        k       p                    �?b�2�tk�?             2@       l       m                   �5@�eP*L��?             &@        ������������������������       �                      @        n       o                 @�pX@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        q       v                    �?����X�?             @       r       u                    >@      �?             @       s       t                 �nc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        w       x                  "&d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        z       �                    B@��T���?)            @R@        {       |                   �<@J�8���?             =@        ������������������������       �                      @        }       ~                 ��I/@�G��l��?             5@        ������������������������       �                     @               �                 0�?D@ҳ�wY;�?	             1@        ������������������������       �                     @        �       �                 �|Y>@���Q��?             $@        ������������������������       �                      @        �       �                   @K@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                   �R@"pc�
�?             F@       �       �                   @J@�T|n�q�?            �E@       �       �                    �?R�}e�.�?             :@        ������������������������       �                     �?        �       �                    �? �o_��?             9@       �       �                 ��#[@�q�q�?             8@       �       �                   �H@R���Q�?             4@       �       �                   �F@�KM�]�?             3@       �       �                 `�iJ@"pc�
�?             &@       �       �                   �E@      �?              @       �       �                   �D@r�q��?             @        ������������������������       �                     �?        �       �                  x#J@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             1@        ������������������������       �                     �?        �       �                   @4@����b�?�            �u@        �       �                   �1@�rF���?'            �K@        �       �                 03�0@�t����?             1@        �       �                   �0@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             "@        �       �                 ��Y @�d�����?             C@       �       �                   �2@�q�q�?             >@        �       �                  s@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �? �o_��?             9@        �       �                 �{@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �3@�GN�z�?             6@       �       �                 �?�@�	j*D�?             *@       ������������������������       �                     @        ������������������������       �և���X�?             @        �       �                 P�@�����H�?             "@        ������������������������       �                     @        �       �                 @3�@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        �                       0��G@̆ꎑ
�?�            @r@       �                          A@���g<�?�            �q@       �       �                   �<@��au���?�            �j@        �       �                    �?���N8�?8             U@        �       �                   �6@"pc�
�?             &@        ������������������������       �                     �?        �       �                 �0@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                     @��pBI�?1            @R@        ������������������������       �        	             (@        �       �                 ���@�]0��<�?(            �N@        �       �                 ���@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �:@�h����?$             L@       ������������������������       �                    �C@        �       �                 pf� @�IєX�?	             1@        ������������������������       �                      @        �       �                   �;@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                     @     |�?R             `@        �       �                   @@@�����H�?             2@       �       �                   �'@�IєX�?             1@        ������������������������       �                     @        �       �                    �?�C��2(�?             &@       �       �                 ��,@�����H�?             "@       �       �                 �|�=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �                        03�5@��2(&�?F            �[@       �       �                 �|Y=@t����?D            �Z@        �       �                    �?      �?             $@        ������������������������       �                     @        �       �                 ���"@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�8��8��?>             X@       �       �                 �?�@㺦���?;            @W@       �       �                 �|�=@ ��WV�?"             J@       �       �                 �Y�@���7�?             F@        �       �                    �?؇���X�?             ,@       �       �                 ���@8�Z$���?             *@        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     >@        ������������������������       �                      @        �       �                 �|�=@,���i�?            �D@       �       �                    �? ��WV�?             :@        ������������������������       �                     @        �       �                 ��) @�nkK�?             7@       ������������������������       �                     *@        �       �                 pf� @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?������?             .@        ������������������������       �                      @        �       �                   �?@�	j*D�?             *@        ������������������������       �                     @        �       �                   @@@ףp=
�?             $@       �       �                 ��I @r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                  S�-@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              03�7@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                  @ �й���?-            @R@                                 �?�g�y��?             ?@                               @D@`2U0*��?             9@        ������������������������       �                     (@              	                `f�)@$�q-�?
             *@        ������������������������       �                     @        
                        �*@�����H�?             "@                                G@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     E@                              p�O@և���X�?             @                              �|�>@      �?             @                             �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������}<����?�/���?br1���?g���Q��?      �?      �?      �?                      �?6eMYS��?���)k��?�������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?�m۶m��?UUUUUU�?�������?      �?                      �?              �?�������?�\V���?)f>���?�L�౼�?�����?������?W�+�Ʌ?��Q�٨�?�q�q�?��8��8�?              �?;�;��?�؉�؉�?              �?      �?      �?      �?                      �?              �?      �?      �?�i��F�?	�=����?      �?      �?�?<<<<<<�?              �?�?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?      �?                      �?              �?��+Q��?�ڕ�]��?              �?^Cy�5�?Cy�5��?R���Q�?���Q��?<<<<<<�?�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ى�؉��?;�;��?�������?�������?�q�q�?9��8���?      �?      �?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?      �?                      �?4և����?������?(������?6��P^C�?�������?�������?      �?                      �?��Moz��?��,d!�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �?�?              �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?        S�-��R�?�Hk���?O��N���?b'vb'v�?��{���?�B!��?              �?���=��?GX�i���?F]t�E�?t�E]t�?�������?333333�?      �?              �?      �?              �?      �?              �?        9��8���?�8��8��?]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?�m۶m��?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �B�
*�?�z��ի�?|a���?�rO#,��?              �?��y��y�?1�0��?      �?        �������?�������?              �?333333�?�������?      �?              �?      �?      �?                      �?/�袋.�?F]t�E�?���)k��?6eMYS��?'vb'vb�?�;�;�?      �?        
ףp=
�?�Q����?�������?�������?333333�?333333�?�k(���?(�����?/�袋.�?F]t�E�?      �?      �?�������?UUUUUU�?      �?        �������?�������?      �?                      �?      �?      �?      �?              �?                      �?              �?      �?              �?                      �?��n^���?����K�?yJ���?�־a��?<<<<<<�?�?      �?      �?              �?      �?              �?        Cy�5��?y�5���?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?
ףp=
�?�Q����?UUUUUU�?UUUUUU�?      �?                      �?�袋.��?]t�E�?vb'vb'�?;�;��?      �?        ۶m۶m�?�$I�$I�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?        *T�P�B�?�^�z��?z�����?/<!W�³?0��>���?~�	�[�?��y��y�?�a�a�?/�袋.�?F]t�E�?              �?�������?�������?      �?                      �?���Ǐ�?����?      �?        \2�h��?;ڼOqɠ?�������?�������?      �?                      �?۶m۶m�?�$I�$I�?      �?        �?�?      �?        �q�q�?�q�q�?              �?      �?             ��?      �?�q�q�?�q�q�?�?�?      �?        ]t�E�?F]t�E�?�q�q�?�q�q�?�������?�������?              �?      �?              �?              �?                      �?��.���?t�E]t�?y+�R�?:�&oe�?      �?      �?              �?�������?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?�]v�e��?EM4�D�?O��N���?;�;��?�.�袋�?F]t�E�?۶m۶m�?�$I�$I�?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?        �����?8��18�?O��N���?;�;��?      �?        �Mozӛ�?d!Y�B�?      �?        �������?�������?              �?      �?        wwwwww�?�?      �?        vb'vb'�?;�;��?              �?�������?�������?�������?UUUUUU�?      �?      �?      �?              �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?              �?      �?        ����Ǐ�?����?��{���?�B!��?���Q��?{�G�z�?      �?        �؉�؉�?;�;��?      �?        �q�q�?�q�q�?�������?�������?UUUUUU�?UUUUUU�?      �?              �?              �?              �?        �$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�	3 hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                 `fK@�3)0�F�?�           8�@              _                 `f�$@4�^��\�?v           x�@                                  �0@^f�(�7�?�            @o@                                   �?�q�q�?             (@       ������������������������       �                     @                                pf�@և���X�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        	       0                 �̌@�?��,�?�            �m@       
                           �?�<ݚ�?S            @]@                                X��B@�+e�X�?             9@                                  �?�q�q�?             8@                                 �2@�㙢�c�?             7@                                P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   8@؇���X�?             5@        ������������������������       �                     "@                                   �?      �?
             (@       ������������������������       �                      @                                �&B@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?               '                 ��@�c:��??             W@              &                    �?P���Q�?5             T@                                   �?������?            �B@                                 �5@      �?             0@        ������������������������       �                      @        ������������������������       �                     ,@                #                 �|Y=@�����?
             5@        !       "                  ��@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        $       %                 03�@�IєX�?             1@        ������������������������       �                      @        ������������������������       ���S�ۿ?             .@        ������������������������       �                    �E@        (       +                 �?$@      �?
             (@        )       *                 �|Y>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ,       -                 P�N@      �?              @        ������������������������       �                     @        .       /                   �>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        1       N                 `�X!@�R����?K            @^@       2       7                 �?�@8v�YeK�?;            �W@        3       6                 �|Y=@P�Lt�<�?             C@        4       5                   �<@�}�+r��?
             3@       ������������������������       �        	             2@        ������������������������       �                     �?        ������������������������       �                     3@        8       9                    �?x�}b~|�?&            �L@        ������������������������       �                      @        :       ;                    �?�C��2(�?$            �K@        ������������������������       �                     �?        <       A                 @3�@h�WH��?#             K@        =       >                    :@      �?              @        ������������������������       �                     @        ?       @                   �?@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        B       C                   �:@�nkK�?             G@        ������������������������       �                     1@        D       E                    <@ 	��p�?             =@        ������������������������       �                     �?        F       M                 �|�=@h�����?             <@        G       H                 �|Y=@�8��8��?	             (@        ������������������������       �                     �?        I       J                 ��) @�C��2(�?             &@       ������������������������       �                      @        K       L                 pf� @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             0@        O       ^                    �?�θ�?             :@       P       Q                  Se!@��+7��?             7@        ������������������������       �                      @        R       S                 ���"@��s����?             5@        ������������������������       �                     @        T       Y                    :@����X�?	             ,@       U       X                    �?�����H�?             "@       V       W                  �#@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        Z       [                    �?���Q��?             @        ������������������������       �                     �?        \       ]                   �?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        `       o                    @�߽���?�            Pu@        a       h                    �?z�G�z�?             >@       b       g                    @ףp=
�?             4@       c       d                 03�=@�}�+r��?             3@       ������������������������       �                     ,@        e       f                 ��T?@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        i       j                    �?���Q��?             $@        ������������������������       �                     @        k       l                 ף�?؇���X�?             @        ������������������������       �                     @        m       n                 ��:@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        p       �                    �?�`���?�            ps@        q       t                    '@     ��?N             `@        r       s                     @�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        u       �                     @z)�J'c�?I            @]@       v       �                   �H@�x
�2�?.            �R@       w       x                   �7@6uH���?)             O@        ������������������������       �                     4@        y       �                  �v7@���H��?             E@       z       �                    �?z�G�z�?             9@       {       |                    �?���N8�?             5@        ������������������������       �                     @        }       ~                   �9@�t����?             1@        ������������������������       �                     �?               �                   @1@      �?             0@       �       �                   �B@8�Z$���?	             *@       ������������������������       �                     $@        �       �                   �*@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        �       �                   �I@      �?             (@        �       �                 03�3@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?v ��?            �E@        �       �                 �|Y=@�q�q�?             "@       �       �                    5@z�G�z�?             @        �       �                 �&�)@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                  S�2@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   @C@j���� �?             A@       �       �                    �?� �	��?             9@        ������������������������       �                     @        �       �                 ���5@�G��l��?             5@        �       �                 �|�<@�	j*D�?             *@        ������������������������       �                     @        ������������������������       �                     "@        �       �                    A@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?hau��?q            �f@        �       �                   �;@�t����?             A@        �       �                    �?      �?              @       �       �                    �?؇���X�?             @       �       �                     @z�G�z�?             @        �       �                 �܅6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     @8�Z$���?             :@       �       �                 p�i@@�8��8��?             8@       �       �                  �>@�t����?	             1@       �       �                    �?      �?             0@       �       �                   �@@@4և���?             ,@       ������������������������       �                     &@        �       �                   �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   @R@h8"J{�?\            �b@       �       �                 ��D:@\�JЂ.�?[            `b@       �       �                    �? ���v��?=            �X@       �       �                    �?H��2�?:            @W@       �       �                    �?���N8�?3             U@        �       �                   `3@�q�q�?             @        ������������������������       �                     �?        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�=@ 7���B�?0            @T@        �       �                   �+@Du9iH��?            �E@        �       �                   �(@@�0�!��?
             1@        �       �                   �2@      �?              @        ������������������������       �                     @        �       �                   �5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y<@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     :@        ������������������������       �                     C@        ������������������������       �                     "@        �       �                 �̌4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             H@        ������������������������       �                     �?        �       �                   �>@�*/�8V�?            �G@        �       �                    K@ҳ�wY;�?             1@       �       �                     �?d}h���?	             ,@       ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     @        �       �                     �?(;L]n�?             >@       �       �                 �|�<@ ��WV�?             :@        �       �                 `f�D@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?E             ^@       �       �                 �|�=@�\=lf�?&            �P@        �       �                 �|�:@�g�y��?             ?@       ������������������������       �        
             4@        �       �                      @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     B@        �                           �?��k��?            �J@       �                         �H@X��ʑ��?            �E@       �       
                   �?���|���?            �@@       �                          �?���Q��?             >@       �       �                  �}S@      �?             8@        �       �                    >@�C��2(�?             &@        �       �                 Ј�Q@z�G�z�?             @       �       �                 0��N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �                       p�w@�n_Y�K�?             *@       �       �                   �8@���!pc�?             &@        ������������������������       �                     @                                 �D@      �?             @                                �?      �?             @                             Ȫ�c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @              	                �̾w@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@                                �7@�z�G��?             $@        ������������������������       �                     @                                 �?      �?             @                             �|�;@���Q��?             @        ������������������������       �                      @                              �|�>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������Rl���?�[�'��?e
�d�?5���7��?�&1��?Zd;�O��?UUUUUU�?UUUUUU�?              �?�$I�$I�?۶m۶m�?      �?              �?      �?����?��o��o�?9��8���?�q�q�?���Q��?R���Q�?�������?UUUUUU�?d!Y�B�?�7��Mo�?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?      �?      �?                      �?      �?              �?        Y�B���?8��Moz�?ffffff�?�������?��g�`��?к����?      �?      �?              �?      �?        =��<���?�a�a�?      �?      �?      �?                      �?�?�?      �?        �������?�?      �?              �?      �?      �?      �?              �?      �?              �?      �?      �?        �������?�������?      �?                      �?�������?���!pc�?��sK���?�a�+�?���k(�?(�����?�5��P�?(�����?      �?                      �?      �?        �YLg1�?Lg1��t�?      �?        ]t�E�?F]t�E�?      �?        ��^B{	�?B{	�%��?      �?      �?      �?        �������?333333�?              �?      �?        �Mozӛ�?d!Y�B�?      �?        ������?�{a���?              �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?        ]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ى�؉��?�؉�؉�?zӛ����?Y�B��?              �?z��y���?�a�a�?      �?        �m۶m��?�$I�$I�?�q�q�?�q�q�?�������?�������?      �?                      �?      �?        �������?333333�?      �?              �?      �?              �?      �?              �?        %�L2�$�?��f�m��?�������?�������?�������?�������?(�����?�5��P�?              �?�������?�������?      �?                      �?      �?        �������?333333�?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        �ںK|_�?J�hA�?      �?      �?]t�E�?F]t�E�?              �?      �?        �)��)��?7k�6k��?o0E>��?�n0E>�?��RJ)��?k���Zk�?              �?��y��y�?�0�0�?�������?�������?��y��y�?�a�a�?              �?�������?�������?      �?              �?      �?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?        G�w��?qG�w��?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?�������?ZZZZZZ�?)\���(�?�Q����?              �?1�0��?��y��y�?;�;��?vb'vb'�?      �?                      �?      �?      �?      �?                      �?      �?        ��o���?��Y@�H�?�������?�������?      �?      �?�$I�$I�?۶m۶m�?�������?�������?      �?      �?      �?                      �?              �?              �?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?<<<<<<�?�?      �?      �?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?                      �?Y���a��?���DxR�?W�7�L�?gG-B���?�y;Cb�?1ogH�۩?�~�駟�?X`��?��y��y�?�a�a�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        	�%����?h/�����?qG�w��?w�qGܱ?ZZZZZZ�?�������?      �?      �?      �?              �?      �?              �?      �?        9��8���?�q�q�?      �?                      �?      �?              �?              �?        �������?UUUUUU�?              �?      �?              �?      �?      �?        �٨�l��?AL� &W�?�������?�������?۶m۶m�?I�$I�$�?              �?      �?              �?        �������?�?O��N���?;�;��?�������?UUUUUU�?              �?      �?              �?              �?                      �?      �?      �?g��1��?"=P9���?�B!��?��{���?              �?F]t�E�?]t�E�?              �?      �?                      �?oe�Cj��?"5�x+��?�}A_�?��}A�?F]t�E�?]t�E]�?�������?333333�?      �?      �?F]t�E�?]t�E�?�������?�������?      �?      �?              �?      �?                      �?              �?;�;��?ى�؉��?F]t�E�?t�E]t�?      �?              �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?      �?      �?      �?                      �?              �?      �?        ffffff�?333333�?      �?              �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       :                     �?�_%����?�           8�@                                   �?Bԅ���?s            �g@                                 "�b@x��B�R�?7            �V@                                  �?@	tbA@�?+            @Q@                                03�=@h�����?             <@        ������������������������       �                     �?        ������������������������       �                     ;@        ������������������������       �                    �D@        	       
                    $@�C��2(�?             6@        ������������������������       �                      @        ������������������������       �                     4@               7                    �?X&$�E�?<            �X@                               `fF:@f���M�?9            @W@        ������������������������       �                     $@               2                    �?�)��V��?4            �T@                                  �?X�<ݚ�?,             R@                                   N@�n_Y�K�?             :@                               �D�G@8����?             7@                                 Y>@���Q��?             $@        ������������������������       �                     @                                   C@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  �5@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @               '                  i?@�LQ�1	�?             G@               "                   @=@�q�q�?
             2@               !                 `f�;@X�<ݚ�?             "@                                   J@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        #       &                 �|Y=@�����H�?             "@        $       %                    <@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        (       -                 ��9L@؇���X�?             <@       )       ,                 �|�<@���}<S�?             7@        *       +                 `f�D@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@        .       1                    C@���Q��?             @       /       0                    >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        3       6                    �?�C��2(�?             &@       4       5                    >@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        8       9                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ;       �                  �#@��+�<�?S           H�@        <       W                    �?�����?�            �k@        =       F                   �7@�0u��A�?)             N@        >       E                    �?�<ݚ�?             "@       ?       B                    �?�q�q�?             @        @       A                 ��y@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        C       D                 ��}@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        G       L                    �?�\�u��?#            �I@        H       I                 ���@��S�ۿ?
             .@        ������������������������       �                     @        J       K                    �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        M       R                 03s@�X�<ݺ?             B@       N       Q                 �|Y=@      �?             @@        O       P                   �<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     <@        S       V                 ��� @      �?             @       T       U                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        X       c                    �?؇���X�?r             d@        Y       b                    �?���Q��?             4@       Z       [                  s@�t����?             1@        ������������������������       �                     @        \       a                 �|Y>@؇���X�?             ,@       ]       `                 ���@$�q-�?             *@        ^       _                 �|Y9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             $@        ������������������������       �                     �?        ������������������������       �                     @        d       k                 �?�@�*/�8V�?b            �a@       e       j                   �8@�(�Tw�?9            �S@        f       i                 ���@ �q�q�?             8@        g       h                 �&b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �        $             K@        l       s                   �4@�<ݚ�?)            �O@        m       r                 ��Y @      �?             0@        n       o                   �2@؇���X�?             @        ������������������������       �                     @        p       q                 @3�@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        t       {                 ��) @t/*�?            �G@       u       z                   �B@���}<S�?             7@       v       w                   �>@���7�?             6@       ������������������������       �        
             ,@        x       y                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        |       }                 �|Y=@      �?             8@        ������������������������       �                     "@        ~       �                   �?@���Q��?             .@               �                 �|�=@���Q��?             $@       �       �                 pf� @և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?Fx$(�?�            �r@        �       �                     @�f7�z�?Z             b@        �       �                    6@�r����?(             N@       �       �                   �J@�<ݚ�?             B@       �       �                 `f�)@@�0�!��?             A@        ������������������������       �                     .@        �       �                   @4@�����?             3@       �       �                   �*@�E��ӭ�?             2@       �       �                    �?�n_Y�K�?             *@       �       �                    ;@�eP*L��?             &@        ������������������������       �                     @        �       �                   �A@      �?              @       ������������������������       �                     @        �       �                    D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        �       �                    @Ї?��f�?2            @U@        �       �                    �?r�q��?             (@        ������������������������       �                     @        �       �                    �?      �?              @        �       �                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 `f�:@z�G�z�?             @        ������������������������       �                      @        �       �                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?X~�pX��?*            @R@        �       �                 �|�;@�P�*�?             ?@        �       �                 �&�)@      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        �       �                    .@���y4F�?             3@        �       �                 ���*@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ��1@�r����?	             .@       ������������������������       �                     $@        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 ���4@���H��?             E@        �       �                   �;@������?             .@        �       �                   �0@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|Y>@ףp=
�?             $@       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 X��@@ 7���B�?             ;@       ������������������������       �        
             0@        �       �                    @�C��2(�?             &@        ������������������������       �                     @        �       �                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @�~R��w�?^            `c@        �       �                    �?��2(&�?             6@       �       �                   �C@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        �       �                 p��D@�<ݚ�?             "@       �       �                    @      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @`�bV��?R            �`@       �       �                    &@P�Lt�<�?-             S@        �       �                    5@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 �|�=@ ����?%            @P@        �       �                    �? 7���B�?             ;@        ������������������������       �                     @        �       �                   �3@���N8�?             5@       �       �                 �|Y<@��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     C@        �       �                    �?Ԫ2��?%            �L@        �       �                 м;4@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                   @@@`�H�/��?"            �I@       �       �                    �?��hJ,�?             A@       �       �                    �?8�Z$���?             :@       �       �                    �?�S����?             3@        �       �                   `3@z�G�z�?             @        ������������������������       �                     @        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �T�C@؇���X�?
             ,@       ������������������������       �                     (@        ������������������������       �                      @        �       �                 `f2@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    #@      �?              @        �       �                 83�@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             1@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������z���� �?@Bx��?�X�0Ҏ�?�S��8�?��?�����?ہ�v`��?�%~F��?�$I�$I�?�m۶m��?      �?                      �?              �?F]t�E�?]t�E�?      �?                      �?b�ΐ���?;Cb�ΐ�?��RJ)��?��Zk���?      �?        ]V��F�?GS��r�?r�q��?�q�q�?ى�؉��?;�;��?8��Moz�?d!Y�B�?333333�?�������?              �?۶m۶m�?�$I�$I�?      �?                      �?;�;��?�؉�؉�?      �?                      �?      �?        Nozӛ��?d!Y�B�?UUUUUU�?UUUUUU�?r�q��?�q�q�?۶m۶m�?�$I�$I�?              �?      �?              �?        �q�q�?�q�q�?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?ӛ���7�?d!Y�B�?333333�?�������?              �?      �?              �?        333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ]t�E�?F]t�E�?۶m۶m�?�$I�$I�?              �?      �?              �?        UUUUUU�?�������?      �?                      �?6��8,�?�� ���?��V��V�?}�}��?�������?�������?�q�q�?9��8���?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?      �?                      �?              �?�������?�?�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        ��8��8�?�q�q�?      �?      �?      �?      �?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        ۶m۶m�?�$I�$I�?333333�?�������?�������?�������?              �?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?r1����?m�w6�;�?p��o���?�A�A�?�������?UUUUUU�?      �?      �?      �?                      �?      �?              �?        9��8���?�q�q�?      �?      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?              �?        �;����?W�+���?ӛ���7�?d!Y�B�?�.�袋�?F]t�E�?      �?              �?      �?              �?      �?                      �?      �?      �?      �?        333333�?�������?�������?333333�?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?        ףp=
��?R���Q�?a���{�?O#,�4��?�?�������?�q�q�?9��8���?�������?ZZZZZZ�?              �?^Cy�5�?Q^Cy��?r�q��?�q�q�?ى�؉��?;�;��?]t�E�?t�E]t�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?              �?                      �?�������?�������?UUUUUU�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�^�z���?�B�
*�?�Zk����?�RJ)���?      �?      �?              �?      �?        (������?6��P^C�?      �?      �?              �?      �?        �?�������?              �?�������?333333�?              �?      �?        �0�0�?��y��y�?wwwwww�?�?�������?333333�?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?	�%����?h/�����?      �?        ]t�E�?F]t�E�?      �?              �?      �?              �?      �?        �4�M�?�,���?t�E]t�?��.���?;�;��?�؉�؉�?              �?      �?        �q�q�?9��8���?      �?      �?              �?      �?              �?        ��f��?�3�τ?�?���k(�?(�����?]t�E�?F]t�E�?              �?      �?         �����? �����?	�%����?h/�����?      �?        ��y��y�?�a�a�?�������?�?      �?                      �?      �?              �?        $���>��?p�}��?      �?      �?              �?      �?        �������?�?KKKKKK�?�������?;�;��?;�;��?(������?^Cy�5�?�������?�������?      �?              �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?              �?      �?      �?      �?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��~hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                  x#J@�C��ӽ�?�           8�@              ;                 ���"@�P�2�?i           P�@                                   �?�.�PI�?�            �m@                                   �?�z�G��?             D@       ������������������������       �                     8@                                �|Y>@      �?
             0@                                  ;@z�G�z�?	             .@                                 �9@�z�G��?             $@       	       
                 pf�@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               $                 ��]@l}N+V5�?�            �h@                               �|Y=@���N8�?E            @Z@                                ���@�����?             E@        ������������������������       �        	             ,@                                  �<@؇���X�?             <@                               ��@�����H�?             ;@        ������������������������       �                     �?                                  �6@$�q-�?             :@                                   �?r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     ,@        ������������������������       �                     �?               #                 �|�=@ ������?*            �O@                                  �? qP��B�?            �E@       ������������������������       �                     7@                                     @P���Q�?             4@       ������������������������       �                     &@        !       "                 ��,@�����H�?             "@       ������������������������       �                     @        ������������������������       �z�G�z�?             @        ������������������������       �                     4@        %       8                 @3�@Ʋ(>^�?;            @W@       &       )                    �?�T`�[k�?!            �J@        '       (                 �|Y=@      �?             (@        ������������������������       �                     @        ������������������������       �                     @        *       1                 �?�@�p ��?            �D@       +       0                   �@(;L]n�?             >@        ,       /                    �?      �?              @       -       .                    >@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     6@        2       5                    :@�eP*L��?             &@        3       4                   �4@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        6       7                   �?@      �?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        9       :                    �?P���Q�?             D@       ������������������������       �                     C@        ������������������������       �                      @        <       y                    �?�q�q�?�            �u@        =       R                     @*(�"u9�?^             c@       >       O                    L@ ,U,?��?0            �T@       ?       B                    �?H�!b	�?.            @T@        @       A                   �H@@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        C       N                    �?�����?%            �P@       D       E                    �?$�q-�?            �C@        ������������������������       �                      @        F       G                     �?�L���?            �B@        ������������������������       �                     @        H       M                   �;@�C��2(�?            �@@        I       L                   �7@���!pc�?             &@       J       K                   �'@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     6@        ������������������������       �                     <@        P       Q                   �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       t                  ��8@B� ��?.            �Q@       T       s                    @��WV��?"             J@       U       `                    �?��e�B��?!            �I@        V       [                    �?@�0�!��?             1@       W       Z                  S�-@      �?              @        X       Y                 ���,@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        \       _                 `�@1@�<ݚ�?             "@        ]       ^                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        a       j                 �|Y=@j���� �?             A@       b       i                   @1@��<b���?             7@       c       h                 pff0@     ��?             0@       d       g                   �*@d}h���?             ,@       e       f                   �3@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        k       r                   @B@"pc�
�?             &@       l       m                   �>@ףp=
�?             $@        ������������������������       �                     @        n       q                    �?r�q��?             @       o       p                 03�1@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        u       v                 ��T?@�����H�?             2@       ������������������������       �                     $@        w       x                 ��p@@      �?              @        ������������������������       �                      @        ������������������������       �                     @        z       �                    @�����D�?s            `h@        {       |                    �?�E��ӭ�?
             2@        ������������������������       �                     �?        }       ~                     @�t����?	             1@        ������������������������       �                     @               �                    @�n_Y�K�?             *@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                 pf�@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     @        �       �                 ��T?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    $@L(ݧa��?i             f@        �       �                   �<@      �?             (@        ������������������������       �                     @        �       �                   �?@�q�q�?             "@       �       �                 �|�=@؇���X�?             @       �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 �D B@�Uk���?c            �d@       �       �                   �R@ Ϸ�~�?V             b@       �       �                    �?h��@D��?U            �a@        �       �                     @�c�Α�?             =@       �       �                 �|�=@R���Q�?             4@       �       �                 �ܵ<@�z�G��?             $@       ������������������������       �                     @        �       �                 ��2>@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    '@X�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?����X�?             @       �       �                 �&�)@�q�q�?             @        ������������������������       �                      @        �       �                 �0@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?ЮN
��?D            @\@        �       �                    �?؇���X�?             @       �       �                 X��E@�q�q�?             @       �       �                   `3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @A@����??            �Z@       �       �                    )@��FM ò?>            @Z@        ������������������������       �                     �?        �       �                 ��D:@��9J���?=             Z@       �       �                   �*@��'�`�?1            �T@        �       �                 �|�=@�?�|�?            �B@        �       �                    �?@4և���?
             ,@       �       �                   �(@$�q-�?	             *@        ������������������������       �                     @        �       �                 �|�<@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                     G@        �       �                     �?�����?             5@       �       �                   @K@r�q��?             (@       �       �                   `G@      �?              @       �       �                 X�,@@؇���X�?             @        ������������������������       �                     @        �       �                    D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        �       �                 ��!T@2]��a�?P            @_@        �       �                 `��M@���@M^�?'             O@        �       �                   �4@PN��T'�?             ;@        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�C��2(�?             6@        ������������������������       �                     (@        �       �                    �?z�G�z�?             $@        ������������������������       �                     �?        �       �                      @�<ݚ�?             "@       �       �                 `�iJ@z�G�z�?             @        ������������������������       �                     �?        �       �                 `f�K@      �?             @       �       �                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�>@      �?             @       �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?և���X�?            �A@        �       �                 0�S@������?             1@       �       �                    �?�8��8��?	             (@       ������������������������       �                     "@        �       �                   �B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|�:@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �7@�����H�?             2@        ������������������������       �                     @        �       �                    �?r�q��?	             (@        �       �                 ���Q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�? Da�?)            �O@       �       �                    �?�Ń��̧?             E@        ������������������������       �                     4@        �       �                 ���a@���7�?             6@       ������������������������       �                     ,@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �                       03c@�q�q�?             5@       �                         @G@8�Z$���?             *@       �                          �?      �?              @                              Ј�V@���Q��?             @        ������������������������       �                     �?                                �5@      �?             @                             �y[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        	      
                X�,@@      �?              @        ������������������������       �                     @                                �B@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub���������������sI,�?��m��?슍���?(���"��?�@��@��?��F��F�?333333�?ffffff�?              �?      �?      �?�������?�������?ffffff�?333333�?9��8���?�q�q�?              �?      �?                      �?      �?                      �?��3$���?;Cb�ΐ�?��y��y�?�a�a�?=��<���?�a�a�?      �?        ۶m۶m�?�$I�$I�?�q�q�?�q�q�?              �?�؉�؉�?;�;��?�������?UUUUUU�?              �?      �?              �?                      �?��}��}�?AA�?��}A�?�}A_З?      �?        ffffff�?�������?      �?        �q�q�?�q�q�?      �?        �������?�������?      �?        /���.�?EM4�D�?���!5��?"5�x+��?      �?      �?              �?      �?        Q��+Q�?��+Q��?�������?�?      �?      �?�������?�������?      �?                      �?      �?              �?        t�E]t�?]t�E�?333333�?�������?      �?      �?      �?              �?      �?              �?333333�?�������?ffffff�?�������?      �?                      �?�������?�������?�g�g�?w!�v!��?��FS�׮?��ˊ��?�����H�?b�2�tk�?�$I�$I�?n۶m۶�?              �?      �?        ���@��?g��1��?;�;��?�؉�؉�?              �?L�Ϻ��?}���g�?              �?F]t�E�?]t�E�?t�E]t�?F]t�E�?333333�?�������?              �?      �?                      �?              �?              �?      �?      �?      �?                      �?B�A��?|�W|�W�?��N��N�?��؉���?�������?�������?�������?ZZZZZZ�?      �?      �?      �?      �?              �?      �?                      �?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?ZZZZZZ�?��,d!�?��Moz��?      �?      �?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        F]t�E�?/�袋.�?�������?�������?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?                      �?�q�q�?�q�q�?      �?              �?      �?              �?      �?        z�z��?z�z��?r�q��?�q�q�?              �?�������?�������?              �?ى�؉��?;�;��?�������?�������?      �?              �?      �?              �?      �?              �?      �?              �?      �?      �?      �?                      �?�C!����?�z���?      �?      �?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?        ��?����?`�1`�?����?�?8���?��V��?�'�K=�?5�rO#,�?�{a���?333333�?333333�?ffffff�?333333�?      �?        �������?333333�?              �?      �?              �?        �q�q�?r�q��?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?m���M�?4��A�/�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        ��`��}�?�V�9�&�?��~���?8�8��?              �?;�;��?�؉�؉�?1P�M��?��k���?*�Y7�"�?к����?n۶m۶�?�$I�$I�?�؉�؉�?;�;��?      �?        �q�q�?�q�q�?      �?                      �?      �?              �?              �?        =��<���?�a�a�?�������?UUUUUU�?      �?      �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?                      �?      �?              �?                      �?              �?      �?        ����Mb�?+����?�c�1��?�s�9��?h/�����?&���^B�?�������?333333�?              �?      �?        F]t�E�?]t�E�?              �?�������?�������?              �?�q�q�?9��8���?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?�$I�$I�?۶m۶m�?�?xxxxxx�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?      �?                      �?�q�q�?�q�q�?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        AA�?�������?�a�a�?��<��<�?              �?F]t�E�?�.�袋�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?;�;��?;�;��?      �?      �?�������?333333�?      �?              �?      �?      �?      �?      �?                      �?              �?              �?              �?      �?      �?      �?        �������?333333�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                   �R@>AU`�z�?�           8�@                                  @$5;Uʹ�?�            �@                                  �C@���N8�?             E@                               @3�4@r�q��?             B@        ������������������������       �        	             ,@                                   �?���!pc�?             6@        ������������������������       �                     @               	                     @ҳ�wY;�?             1@        ������������������������       �                      @        
                        ��T?@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                   '@pTV�h�?�           Ђ@        ������������������������       �                     2@               g                     @@�F���?~           @�@               ,                    �?���`V8�?�            �m@               +                    �?@4և���?:             U@                                  �?���C��?&            �J@        ������������������������       �        
             (@                                  �;@�p ��?            �D@                                  �6@�z�G��?             $@       ������������������������       �                     @                                  �9@      �?             @                                 �3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?               "                   �'@��a�n`�?             ?@                !                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        #       $                   �B@ 	��p�?             =@        ������������������������       �        	             *@        %       &                   @C@      �?
             0@        ������������������������       �                     �?        '       *                   @F@��S�ۿ?	             .@        (       )                    E@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     ?@        -       f                   �R@(Q��w��?c             c@       .       ?                 ��D:@��)�c{�?b             c@       /       0                     �?�zvܰ?6             V@        ������������������������       �                     "@        1       4                    &@(�5�f��?0            �S@        2       3                    5@�����?             5@        ������������������������       ��q�q�?             @        ������������������������       �        
             2@        5       >                    �? _�@�Y�?$             M@       6       =                   �*@0�)AU��?#            �L@       7       8                   �@@Pa�	�?            �@@       ������������������������       �                     5@        9       :                    �?�8��8��?             (@        ������������������������       �                      @        ;       <                   �A@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     8@        ������������������������       �                     �?        @       Q                    �?     ��?,             P@        A       B                 ��";@      �?             8@        ������������������������       �                     �?        C       F                   �;@��<b���?             7@        D       E                     �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        G       P                    �?�KM�]�?             3@       H       O                    H@�r����?
             .@       I       J                 �ܵ<@      �?              @        ������������������������       �                      @        K       N                    B@�q�q�?             @       L       M                 ���=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        R       e                     �?�z�G��?             D@       S       d                    �?�q�q�?             B@       T       [                   �>@^������?            �A@        U       V                 03k:@���!pc�?             &@        ������������������������       �                     @        W       X                 X��B@      �?              @        ������������������������       �                     @        Y       Z                   @J@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        \       a                 ��9L@r�q��?             8@       ]       `                   �B@ףp=
�?             4@        ^       _                 �|�<@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        b       c                 `f�N@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        h       i                 ���@�L�z��?�            �u@        ������������������������       �                     9@        j       �                   @@@�8|^a=�?�             t@       k       �                    �?ؠ���9�?�            Pq@        l       y                    �?�ҿf���?5            �T@        m       t                 �{&@�q�q�?             ;@       n       o                 �|�9@�����H�?             2@        ������������������������       �                     "@        p       q                  ��@�<ݚ�?             "@        ������������������������       �                     �?        r       s                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        u       x                    �?�<ݚ�?             "@       v       w                 pF�-@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        z       �                 03s@X�Cc�?#             L@       {       ~                   �7@д>��C�?             =@        |       }                   �2@      �?             @        ������������������������       �                     @        ������������������������       �                     @               �                    �?���}<S�?             7@        �       �                 �|=@�����H�?             "@        ������������������������       �                      @        �       �                 ���@؇���X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        �       �                  ��@@4և���?             ,@        ������������������������       �                      @        �       �                 �|Y=@�8��8��?	             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?X�<ݚ�?             ;@       �       �                 03�7@      �?             8@       �       �                    �?
;&����?             7@       �       �                 �|Y=@D�n�3�?             3@        �       �                   �;@�8��8��?             (@       �       �                    3@؇���X�?             @        ������������������������       �                     @        �       �                 �0@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   `3@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@�nQ\�?}            @h@        �       �                    �?v���a�?.            @R@        �       �                 ���@�<ݚ�?             "@        ������������������������       �                     @        �       �                 �&B@�q�q�?             @       �       �                    4@���Q��?             @        ������������������������       �                     �?        �       �                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    ?@      �?(             P@       �       �                 ���@�]0��<�?&            �N@        ������������������������       �                     �?        �       �                 �|�<@ �.�?Ƞ?%             N@       ������������������������       �                    �E@        �       �                 �|�=@�IєX�?             1@       �       �                  sW@      �?
             0@        �       �                 pf�@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|�=@
�cՔ��?O            @^@       �       �                   @1@���?��?I            @[@       �       �                 pff0@NP�<��?8            �T@       �       �                    �?l��
I��?7            @T@        �       �                    �?�\��N��?             3@       �       �                   �9@��S���?	             .@       �       �                  �#@�q�q�?             "@       ������������������������       �                     @        �       �                    4@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�;@r�q��?             @        ������������������������       �                     �?        �       �                 pf&(@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �;@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �0@��a�n`�?+             O@        ������������������������       �      �?             @        �       �                 �|Y=@&y�X���?)             M@       �       �                   �:@      �?             F@       �       �                 0S5 @ףp=
�?             >@        �       �                 @3�@      �?	             (@        �       �                   �4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �3@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@        �       �                 pf� @և���X�?             ,@        ������������������������       �                     @        �       �                   �;@���!pc�?             &@        ������������������������       �                     @        �       �                   �<@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                      @        �       �                    �? ��WV�?             :@        ������������������������       �                     $@        �       �                    �?      �?             0@       �       �                    ;@ףp=
�?             $@        �       �                 0��B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �?@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        �       �                    �?`Ӹ����?!            �F@        �       �                   @C@ףp=
�?	             $@        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �C@��?^�k�?            �A@        �       �                 �?�@��S�ۿ?
             .@        ������������������������       �                     @        �       �                   @B@�����H�?             "@        ������������������������       �                     @        �       �                    @r�q��?             @       �       �                 ��	0@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     4@        �                           �?t�U����?-            �P@       �       �                    �?`Ql�R�?            �G@       ������������������������       �                     D@        �       �                 Ъ�c@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @              
                   �?��Q��?             4@             	                 �6f@���!pc�?             &@                                �?z�G�z�?             $@                                �?���Q��?             @                               �5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                 �?X�<ݚ�?             "@                                �?      �?             @                              �̾w@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                             ���u3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?��6�?��2����?��y��y�?�a�a�?UUUUUU�?�������?              �?t�E]t�?F]t�E�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ��O�?�̫�a��?      �?        8p���?�Ǐ?~�?���u�?�����?�$I�$I�?n۶m۶�?"5�x+��?\�琚`�?              �?��+Q��?Q��+Q�?333333�?ffffff�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �c�1Ƹ?�s�9��?      �?      �?              �?      �?        �{a���?������?              �?      �?      �?      �?        �?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�f�f�?�g�g�?Cy�5��?��k(��?颋.���?t�E]t�?      �?        �=Q���?�&��jq�?=��<���?�a�a�?UUUUUU�?UUUUUU�?      �?        #,�4�r�?�{a���?��Gp�?p�}��?|���?|���?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?              �?              �?              �?      �?      �?      �?              �?��,d!�?��Moz��?      �?      �?              �?      �?        �k(���?(�����?�������?�?      �?      �?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?      �?              �?        ffffff�?333333�?UUUUUU�?UUUUUU�?uPuP�?_�_��?t�E]t�?F]t�E�?              �?      �?      �?              �?      �?      �?      �?      �?      �?        �������?UUUUUU�?�������?�������?      �?      �?              �?      �?              �?              �?      �?              �?      �?              �?              �?                      �?re��?�5���?      �?        Q��/�Z�?^����J�?��V�5.�?�@R˔��?S��rY�?Y1P�M�?UUUUUU�?UUUUUU�?�q�q�?�q�q�?              �?�q�q�?9��8���?      �?              �?      �?              �?      �?        9��8���?�q�q�?      �?      �?      �?                      �?      �?        %I�$I��?�m۶m��?a���{�?|a���?      �?      �?      �?                      �?ӛ���7�?d!Y�B�?�q�q�?�q�q�?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �q�q�?r�q��?      �?      �?�Mozӛ�?Y�B��?(������?l(�����?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?      �?              �?      �?      �?                      �?      �?                      �?��W?�?_\����?ٲe˖-�?�4iҤI�?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?�������?333333�?      �?              �?      �?              �?      �?                      �?      �?      �?\2�h��?;ڼOqɠ?              �?wwwwww�?�?      �?        �?�?      �?      �?�������?�������?      �?              �?      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        �GN�z�?"pc�
�?-�M���?N��ش�?%�����?���\V�?Lh/����?h/�����?�5��P�?y�5���?�������?�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?�������?              �?�������?�������?      �?                      �?      �?      �?              �?      �?        �c�1��?�s�9��?      �?      �?��FX��?�i��F�?      �?      �?�������?�������?      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?              �?        ۶m۶m�?�$I�$I�?      �?        t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?      �?                      �?      �?                      �?O��N���?;�;��?      �?              �?      �?�������?�������?      �?      �?      �?                      �?      �?              �?              �?      �?              �?      �?        ?�>��?l�l��?�������?�������?      �?      �?      �?                      �?      �?        _�_��?�A�A�?�������?�?      �?        �q�q�?�q�q�?      �?        �������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?              �?        g��1��?���-�?W�+�ɕ?}g���Q�?              �?�$I�$I�?۶m۶m�?      �?                      �?ffffff�?�������?t�E]t�?F]t�E�?�������?�������?�������?333333�?      �?      �?      �?                      �?      �?                      �?      �?        �q�q�?r�q��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�DhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K兔h2h3h4hph<�h=Kub��������       F                    �?��ϙLq�?�           8�@                                   �?D������?{            `h@                                    @���(`�?3            �U@       ������������������������       �                     K@                                X�,A@r٣����?            �@@                                  �?�n`���?             ?@                                �|Y6@      �?             $@                                  &@�q�q�?             @        	       
                   �@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                      @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                ���@���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                      @               /                   �;@\�f<t�?H             [@               &                   �=@     ��?             @@                                   @��Q��?             4@        ������������������������       �                     �?               %                    �?p�ݯ��?             3@              $                 ؼC1@j���� �?
             1@              !                    �?��S���?	             .@                                  �6@���|���?             &@                                ��y@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        "       #                 ��}@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        '       ,                 �U�X@�q�q�?             (@       (       +                   �8@؇���X�?             @        )       *                 ���Q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        -       .                   �1@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        0       A                    �?h�˹�?3             S@       1       8                  �>@�#-���?.            �Q@       2       3                 `V8@ _�@�Y�?$             M@       ������������������������       �                    �H@        4       7                     �?�����H�?             "@       5       6                 ��";@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        9       @                    �?�q�q�?
             (@       :       ?                 @�pX@      �?	             $@       ;       >                  xCH@      �?              @       <       =                 p�i@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        B       E                     @      �?             @       C       D                 �w�q@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        G       �                    �?BV�(��?G            �@        H       U                     @b�/#w�?n            �d@       I       R                 ��1^@�D�e���?>            @U@       J       Q                    �?�(�Tw�?7            �S@       K       P                  �v7@`���i��?             F@        L       M                   �2@���7�?             6@       ������������������������       �                     4@        N       O                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                     A@        S       T                    !@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        V       w                    �?������?0            �T@       W       X                    @�^���U�?#            �L@        ������������������������       �                     @        Y       v                 ���1@����0�?!             K@       Z       a                   �3@k��9�?            �F@        [       `                   �2@�q�q�?             "@       \       _                 ��!@      �?             @       ]       ^                 P��@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        b       s                    �?*O���?             B@       c       p                 ��Y.@�f7�z�?             =@       d       k                 P�@���!pc�?             6@        e       f                 pff@      �?              @        ������������������������       �                      @        g       h                   �7@r�q��?             @        ������������������������       �                     @        i       j                   �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       m                 ��&@@4և���?
             ,@       ������������������������       �                     &@        n       o                 ���*@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        q       r                 �|�;@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        t       u                   �;@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        x       }                    @HP�s��?             9@       y       |                    @�}�+r��?
             3@        z       {                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        ~       �                    @r�q��?             @              �                 ���A@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��P�sK�?�            �u@       �       �                     �?��cˣ��?�            �r@        �       �                 ��9L@P�~D&�?&            �P@       �       �                    R@d��0u��?"             N@       �       �                   �J@$gv&��?!            �M@       �       �                   �>@��+7��?             G@       �       �                   �G@��>4և�?             <@       �       �                 03:@�q�q�?             8@        ������������������������       �                     &@        �       �                   @=@��
ц��?	             *@       �       �                    D@���Q��?             $@       �       �                 03k:@      �?             @        ������������������������       �                     �?        �       �                 �|�<@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �F@r�q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `fFJ@�X�<ݺ?             2@       ������������������������       �                     (@        �       �                   @K@r�q��?             @       �       �                    7@�q�q�?             @        ������������������������       �                     �?        �       �                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     �?        �       �                 �|Y>@����X�?             @        ������������������������       �                     �?        �       �                 ���R@r�q��?             @       �       �                 03�M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @��xJ_�?�             m@        �       �                    4@ܷ��?��?$             M@        �       �                   �2@�z�G��?             $@       ������������������������       �                     @        ������������������������       �      �?             @        �       �                   @D@      �?             H@       ������������������������       �                     >@        �       �                   �*@r�q��?             2@       �       �                    G@���!pc�?             &@        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �2@ >�֕�?o            �e@        �       �                 ��@�z�G��?             $@        ������������������������       �                     @        �       �                 ��Y @      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�=@�ۊ�̴?g            �d@       �       �                   �;@��7�K¨?K            @^@       �       �                 ���@�nkK�?,            @Q@        �       �                 ���@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �:@�g�y��?&             O@       �       �                 @3�@��v$���?%            �N@       ������������������������       �                    �A@        �       �                 0S5 @ ��WV�?             :@        �       �                   �4@�8��8��?             (@        ������������������������       �      �?              @        ������������������������       �                     $@        ������������������������       �        
             ,@        ������������������������       �                     �?        ������������������������       �                     J@        �       �                 �?�@�C��2(�?             F@        ������������������������       �                     4@        �       �                   @@@r�q��?             8@        �       �                   �?@և���X�?             @        ������������������������       �                      @        ������������������������       ����Q��?             @        ������������������������       �                     1@        �       �                    @ \� ���?             �H@       �       �                 `��S@��+7��?             G@       �       �                    #@��s����?             E@        �       �                    @�q�q�?
             (@        �       �                 �G�?���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @       �       �                 ���7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��9B@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     >@        ������������������������       �                     @        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������Ӭ����?�X�>��?_�^��?�����?Ȥx�L��?g��o��?              �?|���?>���>�?�c�1��?�9�s��?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?        �a�a�?��y��y�?      �?                      �?      �?        ��Kh/�?&���^B�?      �?      �?�������?ffffff�?      �?        ^Cy�5�?Cy�5��?�������?ZZZZZZ�?�?�������?]t�E]�?F]t�E�?�������?�������?      �?                      �?      �?              �?      �?      �?                      �?      �?              �?        �������?�������?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?              �?      �?        ^Cy�5�?�5��P�?�A�A�?_�_�?#,�4�r�?�{a���?      �?        �q�q�?�q�q�?�������?UUUUUU�?              �?      �?              �?        �������?�������?      �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?              �?              �?      �?333333�?�������?      �?                      �?              �?�/����?��/���?E���w��?^�/7Ā�?�???????�?�A�A�?p��o���?F]t�E�?F]t�E�?F]t�E�?�.�袋�?              �?      �?      �?      �?                      �?              �?              �?�$I�$I�?۶m۶m�?      �?                      �?�v%jW��?��+Q��?c:��,��?:��,���?              �?�Kh/���?Lh/����?�'}�'}�?[�[��?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?                      �?              �?�q�q�?�q�q�?O#,�4��?a���{�?F]t�E�?t�E]t�?      �?      �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?              �?        q=
ףp�?{�G�z�?�5��P�?(�����?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?UUUUUU�?�������?�������?              �?      �?              �?        j0֌@��?Y>�����?`,�Œ_�?�6�i�?kL�*g�?*g��1�?�?�������?[4��}�?��/���?zӛ����?Y�B��?۶m۶m�?I�$I�$�?�������?�������?      �?        �؉�؉�?�;�;�?333333�?�������?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?��8��8�?�q�q�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?                      �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?�k�u��?����S��?��=���?a���{�?ffffff�?333333�?      �?              �?      �?      �?      �?      �?        �������?UUUUUU�?F]t�E�?t�E]t�?�������?333333�?      �?              �?        ��+��+�?�A�A�?ffffff�?333333�?      �?              �?      �?              �?      �?        �^G�u��?��[���?�0�~�4�?���!pc�?�Mozӛ�?d!Y�B�?۶m۶m�?�$I�$I�?      �?                      �?��{���?�B!��?.�u�y�?;ڼOqɐ?      �?        O��N���?;�;��?UUUUUU�?UUUUUU�?      �?      �?      �?              �?                      �?      �?        ]t�E�?F]t�E�?      �?        �������?UUUUUU�?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?        
^N��)�?և���X�?zӛ����?Y�B��?z��y���?�a�a�?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���MhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       R                    �?*�Ⱦ��?�           8�@               9                    �?\_D�
��?�            0p@                                   @�ʥ0�?            �i@                                 �K@�â��,�?K             _@                                  �?p�,�V��?I            @^@        ������������������������       �                     F@                                  �E@�g<a�?1            @S@                                 �;@ ��PUp�?+            �Q@        	                           �? �q�q�?             8@       
                          �7@�IєX�?             1@                                  �/@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                    �G@                                  @F@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               6                 ���1@:~=�P�?4            @T@                                  �?\�CX�?-            �Q@                                  �-@�g�y��?             ?@                                   �?r�q��?             @                                 �,@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     9@                3                    �?      �?             D@       !       *                   �@j���� �?             A@        "       )                 �|�;@      �?	             0@       #       $                 pf�@$�q-�?             *@        ������������������������       �                     @        %       (                 �&B@؇���X�?             @        &       '                    4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        +       .                 ��&@X�<ݚ�?             2@       ,       -                    3@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        /       2                 �|�;@�<ݚ�?             "@        0       1                 @3�,@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        4       5                    <@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        7       8                    �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        :       A                     @X�<ݚ�?#             K@        ;       @                     �?$�q-�?             :@        <       =                    �?r�q��?             (@        ������������������������       �                     @        >       ?                    %@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             ,@        B       G                    �?d}h���?             <@        C       F                    @z�G�z�?             @       D       E                 �|Y=@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        H       Q                    @���}<S�?             7@       I       P                    3@�KM�]�?             3@       J       K                 ��	0@r�q��?             (@        ������������������������       �                     �?        L       M                 ��T?@�C��2(�?             &@       ������������������������       �                     "@        N       O                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        S                          @j̬�b��?$           @|@       T       c                    #@h�!��?!           �{@        U       V                 �Q��?
j*D>�?             :@        ������������������������       �                      @        W       `                    �?      �?             8@       X       [                    @��S���?             .@        Y       Z                     @����X�?             @        ������������������������       �                      @        ������������������������       �                     @        \       ]                    @      �?              @       ������������������������       �                     @        ^       _                 03�6@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        a       b                 ���9@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        d       �                     �?�>4և��?           @z@        e       �                    �?�q�q�?8            @W@       f       q                    �?&:~�Q�?.             S@        g       p                 ��<J@�G�z��?             4@       h       i                 �|�;@d}h���?	             ,@        ������������������������       �                     �?        j       k                 `f&;@8�Z$���?             *@        ������������������������       �                     �?        l       o                    H@�8��8��?             (@       m       n                    C@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        r       s                 ��<:@��X��?"             L@        ������������������������       �                     *@        t       {                   �<@�K��&�?            �E@        u       v                 `f�D@����X�?             @        ������������������������       �                     @        w       x                    7@      �?             @        ������������������������       �                     �?        y       z                   �;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        |       �                   @A@*O���?             B@        }       ~                 �|Y>@�C��2(�?             &@       ������������������������       �                     @               �                   @K@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �D@�q�����?             9@        ������������������������       �                     @        �       �                   �G@8�A�0��?             6@       �       �                   �F@����X�?             ,@        �       �                 ���K@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `f�<@      �?              @       �       �                   �J@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �7@������?
             1@        ������������������������       �                     @        �       �                 �̾w@@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        �       �                     @�	CO���?�            pt@        �       �                    �?��
���?2            �R@       �       �                   �@@��.N"Ҭ?.            @Q@       ������������������������       �                    �C@        �       �                   @A@��S�ۿ?             >@        �       �                    1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �*@ ��WV�?             :@       �       �                   �)@$�q-�?	             *@       ������������������������       �                      @        �       �                    G@z�G�z�?             @        �       �                   @D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     @        �       �                   @@@r�q��?�            �o@       �       �                   �>@����R��?�            `j@       �       �                 �|Y=@0�W���?�            @i@       �       �                    �?�x���_�?L            �]@        �       �                    <@b�2�tk�?             2@       �       �                    �?      �?	             ,@       �       �                   �:@��
ц��?             *@       �       �                   �6@�q�q�?             "@       �       �                    5@z�G�z�?             @       �       �                    0@�q�q�?             @        ������������������������       �                     �?        �       �                 �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �8@      �?             @        ������������������������       �                     �?        �       �                 �0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �<@�:pΈ��?A             Y@       �       �                    �?�KM�]�??            �W@       �       �                 �?�@�Ra����?:             V@        ������������������������       �                    �C@        �       �                 0S5 @�����?             �H@        �       �                 @3�@X�<ݚ�?             2@        �       �                   �4@և���X�?             @        ������������������������       ����Q��?             @        ������������������������       �                      @        �       �                   �4@�eP*L��?             &@       �       �                   �2@      �?              @       �       �                    1@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     @        �       �                   �:@`Jj��?             ?@       ������������������������       �                     :@        �       �                 ��)"@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �̌!@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �? �Cc}�?8             U@       �       �                 �Y5@ףp=
�?5             T@        �       �                 �|�=@@�0�!��?             A@       �       �                 ��@     ��?             @@       �       �                    �?؇���X�?             <@        �       �                 ���@�q�q�?             "@        ������������������������       �                     @        ������������������������       ����Q��?             @        �       �                    �?�}�+r��?             3@       �       �                 ���@      �?             0@        ������������������������       �                     @        ������������������������       �ףp=
�?             $@        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                      @        �       �                 �|�=@�nkK�?             G@       �       �                    �? �#�Ѵ�?            �E@        ������������������������       �                      @        �       �                 ��) @ >�֕�?            �A@       ������������������������       �                     7@        �       �                 �̜!@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �?@�q�q�?             "@        �       �                 pff@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �!B@�q�q�?             @       �       �                 P�@      �?             @        ������������������������       �                     �?        �       �                 pf�'@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        �                          �?������?            �D@       �       �                 �?�@@-�_ .�?            �B@        ������������������������       �                     2@        �                        @3�@�KM�]�?             3@        ������������������������       ��q�q�?             @        ������������������������       �        
             0@        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�����������������?�{d�_�?.�!J��?4�w-F��?|��{�?�{���?�c�1Ƙ?:�s�9�?���k��?ˠT�x�?              �?�cj`?���8+�?��V،?��ۥ���?UUUUUU�?�������?�?�?UUUUUU�?�������?              �?      �?                      �?              �?              �?UUUUUU�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ��E���?�<ݚ�?��V��?=�]���?�B!��?��{���?UUUUUU�?�������?�������?�������?              �?      �?                      �?              �?      �?      �?ZZZZZZ�?�������?      �?      �?;�;��?�؉�؉�?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        r�q��?�q�q�?�q�q�?�q�q�?              �?      �?        �q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?�������?              �?      �?        �������?�������?              �?      �?        �q�q�?r�q��?;�;��?�؉�؉�?UUUUUU�?�������?              �?�q�q�?9��8���?      �?                      �?              �?I�$I�$�?۶m۶m�?�������?�������?      �?      �?              �?      �?                      �?ӛ���7�?d!Y�B�?�k(���?(�����?�������?UUUUUU�?              �?]t�E�?F]t�E�?      �?              �?      �?              �?      �?              �?              �?        ���ZX��?驅��Z�?��4n`��?t�,G~��?b'vb'v�?;�;��?              �?      �?      �?�?�������?�m۶m��?�$I�$I�?              �?      �?              �?      �?              �?      �?      �?              �?      �?        9��8���?�q�q�?              �?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?�k(���?�k(����?�������?�������?I�$I�$�?۶m۶m�?              �?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?                      �?      �?                      �?n۶m۶�?%I�$I��?      �?        ��)kʚ�?���)k��?�$I�$I�?�m۶m��?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?]t�E�?F]t�E�?      �?        �������?�������?      �?                      �?�p=
ף�?���Q��?              �?颋.���?/�袋.�?�m۶m��?�$I�$I�?r�q��?�q�q�?              �?      �?              �?              �?      �?333333�?�������?              �?      �?                      �?xxxxxx�?�?              �?n۶m۶�?�$I�$I�?      �?                      �?��h���?�a\&9�?&�X�%�?O贁N�?�3J���?ہ�v`��?      �?        �������?�?      �?      �?              �?      �?        O��N���?;�;��?�؉�؉�?;�;��?      �?        �������?�������?      �?      �?      �?                      �?      �?              �?              �?        �������?UUUUUU�?��ʣ��?��p�C�?�&��?���g��?�<�"h8�?'u_�?9��8���?�8��8��?      �?      �?�;�;�?�؉�؉�?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?��Q���?�Q����?�k(���?(�����?]t�E]�?]t�E�?      �?        ^N��)x�?����X�?r�q��?�q�q�?�$I�$I�?۶m۶m�?�������?333333�?      �?        t�E]t�?]t�E�?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        ���{��?�B!��?      �?        333333�?�������?              �?      �?              �?        �������?�������?      �?                      �?%I�$I��?۶m۶m�?�������?�������?ZZZZZZ�?�������?      �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        �������?333333�?�5��P�?(�����?      �?      �?      �?        �������?�������?      �?              �?      �?      �?        �Mozӛ�?d!Y�B�?�/����?�}A_Ч?      �?        ��+��+�?�A�A�?      �?        �������?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?p>�cp�?������?S�n0E�?к����?      �?        �k(���?(�����?UUUUUU�?UUUUUU�?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ9M�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       \                    �?\��m͗�?�           8�@               G                    �?03�Z*!�?�            �n@                                   @ʨ����?|             h@                                 �K@ج��w�?G            �\@                                 �B@X'"7��?D             [@       ������������������������       �        1            �T@                                    �?���B���?             :@                                  �?�����H�?             2@        	       
                   �H@      �?              @       ������������������������       �                     @                                   J@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@                                  �3@      �?              @                                 �'@����X�?             @        ������������������������       �                      @                                  �*@���Q��?             @                                  D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                  �L@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                   @����[��?5            �S@        ������������������������       �                     @               *                    �?F�����?1            @R@               %                 �&�)@؇���X�?             <@                                   �?P���Q�?             4@        ������������������������       �                      @        !       "                 �|�9@�X�<ݺ?             2@        ������������������������       �                      @        #       $                 ���@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        &       '                 �|6@      �?              @        ������������������������       �                      @        (       )                  S�-@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        +       D                 �|Y>@��S���?            �F@       ,       -                 ���@Hث3���?            �C@        ������������������������       �                     @        .       ?                   �;@և���X�?            �A@       /       <                   �9@      �?             :@       0       ;                   �6@�q�q�?             2@       1       6                 ��,#@��
ц��?	             *@        2       5                 �&B@      �?              @        3       4                    4@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        7       :                    3@z�G�z�?             @        8       9                 �y�+@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        =       >                 @3�,@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        @       A                   �.@�<ݚ�?             "@       ������������������������       �                     @        B       C                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        E       F                   �A@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        H       M                     @~|z����?$            �J@        I       J                 ���[@�X�<ݺ?             2@       ������������������������       �                     $@        K       L                    $@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        N       S                 �̼6@4�2%ޑ�?            �A@        O       P                 ��Y@���Q��?             $@        ������������������������       �                      @        Q       R                 �|Y=@      �?              @       ������������������������       �                     @        ������������������������       �                      @        T       Y                    @HP�s��?             9@       U       X                 ��p@@���N8�?             5@       V       W                    @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     &@        Z       [                 ���A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ]       l                    @6i��� �?            }@        ^       _                   �5@�q�q�?             2@        ������������������������       �                     @        `       k                  DP@��
ц��?             *@       a       f                    �?�q�q�?             "@        b       e                   �C@���Q��?             @       c       d                   A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        g       j                    @      �?             @       h       i                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        m       �                 ��D:@�6��2��?           �{@       n       �                    �?a�G���?�            �t@        o       �                    �?RB)��.�?            �E@       p       q                     @�ݜ�?            �C@        ������������������������       �                      @        r       w                 ���@$G$n��?            �B@        s       t                 ��y@      �?	             0@        ������������������������       �                     �?        u       v                 �|�9@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        x       �                 �&�)@��s����?             5@       y       �                 83##@      �?	             0@       z       }                 �|Y=@z�G�z�?             .@        {       |                   �<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ~                          @@�C��2(�?             &@        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                     �?�X�<ݺ?�             r@        ������������������������       �                     @        �       �                    �?8�wO�?�            �q@        �       �                     @��S�ۿ?             >@        ������������������������       �                      @        �       �                   `3@@4և���?             <@       ������������������������       �                     :@        ������������������������       �                      @        �       �                   @4@0�!��ú?�            �o@        �       �                 pf� @���5��?"            �L@       �       �                    �?H�V�e��?             A@       �       �                   �2@     ��?             @@        �       �                   �1@���Q��?             $@       �       �                 pf�@؇���X�?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 �?�@��2(&�?             6@       ������������������������       �                     ,@        �       �                   �3@      �?              @        ������������������������       �      �?             @        �       �                 @3�@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     7@        �       �                    �?h�����?~            �h@       �       �                     @�	�(�Z�?x            �g@        �       �                   @@@�NW���?"            �J@        ������������������������       �                     6@        �       �                   �E@��� ��?             ?@       �       �                    1@�<ݚ�?
             2@       �       �                   �'@������?             .@        ������������������������       �                     �?        �       �                   @D@����X�?             ,@       �       �                   �A@z�G�z�?             $@        ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �        	             *@        �       �                 P�N@����?�?V            �`@        ������������������������       �                     F@        �       �                 �Yu@x��B�R�?;            �V@        �       �                    =@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �B@�x�E~�?9            @V@       �       �                 @Q!@����ȫ�?2            �T@       ������������������������       �        %            �N@        �       �                 @3�!@���N8�?             5@        �       �                   �:@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                 @3�@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                      @        �       �                  �>@�e"��?F             ]@        �       �                     �?��J�fj�?            �B@       �       �                    D@�c�Α�?             =@       �       �                   @>@r�q��?
             2@       �       �                 X�,@@�θ�?             *@       �       �                   �<@և���X�?             @        ������������������������       �                     @        �       �                 �ܵ<@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @=@�eP*L��?             &@       �       �                 `f�;@      �?              @       �       �                   �K@      �?             @       �       �                    H@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @I@p`q�q��?0            �S@       �       �                     �?��6}��?'            �N@       �       �                    �?�J��%�?            �H@        �       �                    �?
j*D>�?             :@       �       �                    C@8�A�0��?             6@       �       �                 �|Y<@      �?             0@        �       �                   �8@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �H@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             @        �       �                    B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                  "&d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���R@��<b���?             7@       �       �                   �B@�X�<ݺ?             2@        �       �                 �TaA@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             .@        �       �                 X��@@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �        	             2@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub���������������"`c�?ȃ޺?9�?!�M!�?��~Y��?�P�ݙ��?�+���\�?A�V���?�%��~�?B{	�%��?Lh/����?              �?ى�؉��?��؉���?�q�q�?�q�q�?      �?      �?              �?      �?      �?      �?                      �?              �?      �?      �?�$I�$I�?�m۶m��?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �$I�$I�?۶m۶m�?      �?                      �?5H�4H��?�[��[��?              �?�^�z���?�P�B�
�?�$I�$I�?۶m۶m�?�������?ffffff�?              �?�q�q�?��8��8�?              �?�������?�������?      �?                      �?      �?      �?      �?        UUUUUU�?�������?      �?                      �?�������?�?�i�i�?��-��-�?              �?�$I�$I�?۶m۶m�?      �?      �?UUUUUU�?UUUUUU�?�;�;�?�؉�؉�?      �?      �?333333�?�������?      �?                      �?              �?�������?�������?      �?      �?              �?      �?              �?              �?              �?      �?              �?      �?        9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?      �?        �	�[���?��sHM0�?�q�q�?��8��8�?              �?      �?      �?      �?                      �?�������?�A�A�?�������?333333�?      �?              �?      �?              �?      �?        q=
ףp�?{�G�z�?��y��y�?�a�a�?�������?�������?              �?      �?              �?              �?      �?              �?      �?        �:��S��?_�E�^�?UUUUUU�?UUUUUU�?              �?�؉�؉�?�;�;�?UUUUUU�?UUUUUU�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?      �?      �?                      �?      �?                      �?�Xۿ��?�뜒 ��?Uv�D��?eWMT�U�?S֔5eM�?���)k��?\��[���?�i�i�?      �?        к����?���L�?      �?      �?      �?        �������?�?              �?      �?        z��y���?�a�a�?      �?      �?�������?�������?      �?      �?      �?                      �?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?                      �?��8��8�?�q�q�?      �?        �;�0�?ƿD\n�?�������?�?      �?        n۶m۶�?�$I�$I�?      �?                      �?��0�:�?�����T�?�}��?��Gp�?iiiiii�?ZZZZZZ�?      �?      �?333333�?�������?۶m۶m�?�$I�$I�?      �?              �?      �?              �?��.���?t�E]t�?      �?              �?      �?      �?      �?      �?      �?      �?      �?      �?              �?              �?        �m۶m��?�$I�$I�?������?L� &W�?萚`���?�x+�R�?      �?        �{����?�B!��?9��8���?�q�q�?wwwwww�?�?      �?        �m۶m��?�$I�$I�?�������?�������?�m۶m��?�$I�$I�?      �?              �?      �?      �?              �?        ��I��I�?l�l��?      �?        �����?��?      �?      �?      �?                      �?����G�?p�\��?������?������?      �?        ��y��y�?�a�a�?�������?�������?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?        ������?�FX�i�?к����?�"�u�)�?�{a���?5�rO#,�?UUUUUU�?�������?�؉�؉�?ى�؉��?۶m۶m�?�$I�$I�?              �?      �?      �?      �?              �?      �?              �?      �?                      �?              �?]t�E�?t�E]t�?      �?      �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        
�Z܄�?�3����?�!XG��?;ڼOq��?c}h���?9/����?b'vb'v�?;�;��?颋.���?/�袋.�?      �?      �?r�q��?�q�q�?      �?                      �?      �?        UUUUUU�?�������?              �?      �?              �?      �?      �?      �?              �?      �?              �?      �?              �?      �?        ��,d!�?��Moz��?��8��8�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJpVhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0Kㅔh2h3h4hph<�h=Kub��������       N                 `f�$@�C�"���?�           8�@                                   �?@w��_m�?�            �o@                                  �3@��H�}�?             I@        ������������������������       �                     0@                                  �4@��.k���?             A@        ������������������������       �                     @                                �̌@П[;U��?             =@                                  �?���N8�?             5@       	       
                 ���@������?             1@        ������������������������       �                      @                                03@�r����?
             .@                               �|�9@"pc�
�?             &@        ������������������������       �                      @                                   �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                ���@      �?             @        ������������������������       �                      @                                ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                     @���2j��?�            �i@        ������������������������       �                     �?               9                 �?�@`�a�?�            `i@              ,                    �?�S���?P             ^@               )                    �?      �?             D@               (                   @@R���Q�?             4@              !                   �5@�KM�]�?             3@                                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        "       #                 ���@�IєX�?
             1@        ������������������������       �                      @        $       %                 �|=@�����H�?             "@        ������������������������       �                     @        &       '                 �|�=@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        *       +                 �|Y=@ףp=
�?             4@        ������������������������       �                      @        ������������������������       �                     2@        -       .                    7@�(\����?6             T@        ������������������������       �                     5@        /       2                   �8@���#�İ?&            �M@        0       1                   �@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        3       4                 ��L@�h����?$             L@       ������������������������       �                     ?@        5       8                   �@`2U0*��?             9@        6       7                    >@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     3@        :       ;                    �?b:�&���?2            �T@        ������������������������       �                     @        <       M                   @@@̘SJl��?0            �S@       =       L                 0S%"@j�g�y�?%             O@       >       G                   �>@�I� �?             G@       ?       D                 ��) @      �?             B@       @       C                   �3@���B���?             :@        A       B                   �2@����X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     3@        E       F                   �7@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        H       I                   �?@���Q��?             $@        ������������������������       �                     �?        J       K                 ��I @X�<ݚ�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     1@        O       �                     @�t����?           �|@       P       a                    �?�w��$_�?�            �s@        Q       `                    :@�ㄡ^�?S             a@        R       _                    �?HP�s��?!             I@       S       V                   �2@������?            �D@       T       U                    L@XB���?             =@       ������������������������       �                     <@        ������������������������       �                     �?        W       X                    �?      �?             (@        ������������������������       �                     �?        Y       \                   �7@���!pc�?             &@        Z       [                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ]       ^                   �E@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �        2            �U@        b       u                    ,@hp�ɞ�?m             f@        c       h                    4@�L���?            �B@        d       e                   �2@�q�q�?             @        ������������������������       �                     �?        f       g                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        i       j                   �)@�IєX�?             A@        ������������������������       �        	             (@        k       t                   �*@�C��2(�?             6@       l       m                 �|�<@ףp=
�?             4@        ������������������������       �                     "@        n       o                 �|�=@"pc�
�?             &@        ������������������������       �                     �?        p       q                   �C@ףp=
�?             $@        ������������������������       �                     @        r       s                    G@؇���X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        v       �                    @�I'$;=�?R            �a@       w       �                   �<@4V��X�?Q            `a@        x       �                  "&d@<ݚ)�?             B@       y       �                     �?r٣����?            �@@       z       �                    �?�S����?             3@       {       |                   �8@     ��?	             0@        ������������������������       �                      @        }       ~                   �;@@4և���?             ,@       ������������������������       �                     @               �                 `f�D@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    "@X�Cc�?	             ,@        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?6�"W�u�?;            �Y@       �       �                  x#J@RB)��.�?0            �U@       �       �                  �>@0)RH'�?'            @Q@       �       �                    �?��Q���?             D@        �       �                     �?�����H�?             "@        �       �                 �|�=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   @=@�4�����?             ?@       �       �                 `fF:@      �?             <@        ������������������������       �                     @        �       �                 `f�:@�q�q�?	             5@       �       �                   �K@     ��?             0@       �       �                 X��B@���|���?             &@        ������������������������       �                     @        �       �                   @G@      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     =@        �       �                 �|Y>@j���� �?	             1@        ������������������������       �                     @        �       �                    �?�z�G��?             $@        �       �                 @�pX@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �B@z�G�z�?             @        �       �                    A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                     �?        �       �                    �?$�}�$>�?\            �a@       �       �                 ��Y7@J�����?/            @S@       �       �                   �D@RB)��.�?            �E@       �       �                    �?��s����?             E@       �       �                 P��+@�<ݚ�?             B@        ������������������������       �                      @        �       �                 �|�;@����X�?             <@        �       �                 pff0@�eP*L��?             &@        ������������������������       �                     @        �       �                 ��*4@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                  S�-@�t����?
             1@        ������������������������       �                     �?        �       �                 03�1@      �?	             0@       ������������������������       �                     "@        �       �                    �?؇���X�?             @        �       �                 �|Y>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    @l��\��?             A@        �       �                 ��T?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    A@`Jj��?             ?@       �       �                 �|Y9@h�����?             <@        ������������������������       �                     $@        �       �                    �?�X�<ݺ?             2@        ������������������������       �                     �?        ������������������������       �                     1@        �       �                    @�q�q�?             @        ������������������������       �                     �?        �       �                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?6YE�t�?-            �P@        �       �                 �|Y<@      �?              @       �       �                 �&�)@����X�?             @        ������������������������       �                     �?        �       �                 �0@r�q��?             @        ������������������������       �                     @        �       �                   �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    #@�y��*�?'             M@        �       �                 @3�4@      �?
             0@        ������������������������       �                     @        ������������������������       �                     $@        �       �                 �T�I@�Ń��̧?             E@       ������������������������       �                    �B@        �       �                    ;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������[�e�?���I54�?M&��d2�?�f��l6�?
ףp=
�?{�G�z�?              �?�������?�?      �?        ��=���?�{a���?��y��y�?�a�a�?�?xxxxxx�?      �?        �?�������?F]t�E�?/�袋.�?              �?�q�q�?9��8���?              �?      �?                      �?      �?      �?              �?      �?      �?      �?                      �?      �?        �������?�������?      �?        �^q2��?Ztl��?""""""�?�����ݭ?      �?      �?333333�?333333�?�k(���?(�����?      �?      �?              �?      �?        �?�?      �?        �q�q�?�q�q�?      �?        �������?UUUUUU�?      �?      �?      �?                      �?�������?�������?              �?      �?        333333�?�������?      �?        ��N��?'u_[�?UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?�$I�$I�?      �?        ���Q��?{�G�z�?�������?UUUUUU�?      �?                      �?      �?        �b��7�?o4u~�!�?      �?        �3����?�0���M�?B!�B�?��{���?Y�B���?Nozӛ��?      �?      �?��؉���?ى�؉��?�$I�$I�?�m۶m��?              �?      �?      �?      �?        333333�?�������?      �?                      �?�������?333333�?              �?�q�q�?r�q��?      �?      �?      �?              �?              �?        M?�b�,�?g��:_��?����?r�p7�=�?������?�;�H��?{�G�z�?q=
ףp�?������?�|����?�{a���?GX�i���?              �?      �?              �?      �?              �?t�E]t�?F]t�E�?      �?      �?      �?                      �?�q�q�?9��8���?              �?      �?                      �?              �?�Br��?�z���?}���g�?L�Ϻ��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �?�?      �?        ]t�E�?F]t�E�?�������?�������?      �?        /�袋.�?F]t�E�?              �?�������?�������?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?        ��+��+�?�:��:��?'!����?���n��?�8��8��?��8��8�?|���?>���>�?^Cy�5�?(������?      �?      �?      �?        �$I�$I�?n۶m۶�?              �?�$I�$I�?۶m۶m�?              �?      �?                      �?�m۶m��?%I�$I��?              �?      �?              �?        w��jch�?#>�Tr^�?S֔5eM�?���)k��?��k��?F��Q�g�?333333�?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?        ���Zk��?��RJ)��?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?F]t�E�?]t�E]�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �������?ZZZZZZ�?      �?        333333�?ffffff�?�������?333333�?              �?      �?        �������?�������?      �?      �?              �?      �?                      �?      �?              �?        -)D�{�?���w��?V~B����?S{����?���)k��?S֔5eM�?�a�a�?z��y���?�q�q�?9��8���?              �?�$I�$I�?�m۶m��?t�E]t�?]t�E�?      �?        �$I�$I�?�m۶m��?              �?      �?        �?<<<<<<�?      �?              �?      �?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        ------�?�������?UUUUUU�?UUUUUU�?      �?                      �?���{��?�B!��?�m۶m��?�$I�$I�?      �?        ��8��8�?�q�q�?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        '�l��&�?e�M6�d�?      �?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�4�rO#�?GX�i��?      �?      �?              �?      �?        ��<��<�?�a�a�?      �?        �������?�������?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM%hjh))��}�(h,h/h0M%��h2h3h4hph<�h=Kub������       l                    �?���$ӡ�?�           8�@               !                     @n�8����?�            �n@                                  �?�M8��p�?Y             a@                                ��A@@�E�x�?!            �H@                                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     E@        	                           @����!p�?8             V@        
                            �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                    �? �#�Ѵ�?6            �U@                                   �?�>����?!             K@        ������������������������       �        
             3@                                  �7@(N:!���?            �A@                                 `2@R���Q�?             4@                                 �J@�����H�?             2@                               `f�)@�IєX�?             1@       ������������������������       �                     $@                                  �C@؇���X�?             @                                  �B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                   ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �E@��S�ۿ?	             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     @@        "       ]                    �?8�A�0��?F            �[@       #       0                    �?�P�����?6             U@        $       -                    �?��G���?            �B@       %       &                 �{&@ 	��p�?             =@       ������������������������       �                     3@        '       (                   �-@z�G�z�?             $@        ������������������������       �                     �?        )       *                 �|Y6@�����H�?             "@        ������������������������       �                     @        +       ,                  S�-@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        .       /                    @      �?              @        ������������������������       �                     @        ������������������������       �                     @        1       X                 ���1@֭��F?�?            �G@       2       M                 `f�%@�4F����?            �D@       3       B                   �5@�q�q�?             8@        4       ?                   �4@����X�?             ,@       5       >                   �3@�q�q�?             "@       6       =                    �?      �?              @       7       8                 P��@����X�?             @        ������������������������       �                     @        9       <                   �2@      �?             @       :       ;                 ��!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        @       A                 ��y!@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        C       J                 �?�@���Q��?	             $@       D       E                 ��@z�G�z�?             @        ������������������������       �                      @        F       I                  sW@�q�q�?             @       G       H                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        K       L                  S�"@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        N       U                    �?@�0�!��?	             1@       O       T                   �D@z�G�z�?             $@       P       Q                    /@�����H�?             "@        ������������������������       �                     @        R       S                 �|�;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        V       W                    .@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        Y       Z                    �?r�q��?             @        ������������������������       �                      @        [       \                   �>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ^       a                    �?�θ�?             :@        _       `                 �|Y=@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        b       k                 ��p@@��2(&�?             6@       c       h                    @      �?	             (@       d       g                 ��l4@�����H�?             "@        e       f                 �|�:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        i       j                   @C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        m       �                 ��D:@�����S�?            }@       n       u                    $@�)���?�            u@        o       p                     @؇���X�?             ,@        ������������������������       �                     @        q       t                    @�<ݚ�?             "@        r       s                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        v       �                 �|Y=@x������?�            0t@        w       �                    �?     |�?L             `@        x       {                 ���.@�q�q�?	             (@       y       z                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        |       }                 ؼC1@      �?             @        ������������������������       �                     �?        ~                          �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q3�M��?C             ]@       �       �                     @�:�H:�?@            @[@        �       �                    5@�}�+r��?             3@        �       �                   �2@      �?             @        ������������������������       �                     �?        �       �                   �'@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        �       �                 �?�@�����H�?5            �V@       �       �                   �7@p���?             I@       ������������������������       �                     A@        �       �                   �8@      �?	             0@        �       �                   �@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        �       �                   �0@R���Q�?             D@        ������������������������       �                     �?        �       �                   �:@x�����?            �C@       �       �                 0S5 @\-��p�?             =@        �       �                   �4@      �?	             0@       �       �                 @3�@���Q��?             $@        ������������������������       ��q�q�?             @        �       �                   �3@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             *@        �       �                   �;@���Q��?             $@        ������������������������       �                     @        �       �                 ���"@؇���X�?             @        ������������������������       �                     @        �       �                   �<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��]@࿾��@�?y            `h@        �       �                    �? ��ʻ��?(             Q@        �       �                 ���@@4և���?	             ,@       ������������������������       �                     @        �       �                 �|�=@؇���X�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                      @        ������������������������       �                     K@        �       �                 �|�=@HVĮ���?Q            �_@        �       �                    �?`���i��?             F@       ������������������������       �                    �E@        ������������������������       �                     �?        �       �                   @@@��Lɿ��?8            �T@        �       �                   �@�q�q�?             2@        ������������������������       �                      @        �       �                   �>@      �?             0@        �       �                    �?؇���X�?             @        ������������������������       �                     �?        �       �                     @r�q��?             @        ������������������������       �                      @        �       �                 �̌!@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�q�?             "@       �       �                     @      �?              @        ������������������������       �                      @        �       �                   �?@      �?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     �?        �       �                     @P�2E��?*            @P@       �       �                    �?��?^�k�?            �A@       �       �                   �*@г�wY;�?             A@       �       �                 `f�)@      �?             0@        ������������������������       �                     @        �       �                   �C@�C��2(�?             &@        ������������������������       �                     @        �       �                   �F@؇���X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �        
             2@        ������������������������       �                     �?        �       �                    �?��S�ۿ?             >@        ������������������������       �                     @        �       �                 @3�@HP�s��?             9@        �       �                 �?�@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@        �                           �?PlX=��?P            �_@       �       �                    �?���H.�?;             Y@        �       �                   �:@�����?             C@        �       �                    �?���|���?             &@       �       �                   �8@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @F@�+$�jP�?             ;@       �       �                 p�w@�t����?
             1@       �       �                    C@      �?	             0@       �       �                 �|�=@؇���X�?             ,@       �       �                 ��2>@"pc�
�?             &@        ������������������������       �                     �?        �       �                 �|Y<@ףp=
�?             $@        �       �                 Ъb@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �                          @�g�y��?#             O@       �       �                    @@      �?"             N@        �       �                 `fF<@�q�q�?             8@       �       �                   �J@�t����?
             1@       �       �                 03k:@؇���X�?             ,@        ������������������������       �                     �?        �       �                   �C@8�Z$���?             *@        ������������������������       �                     @        �       �                   @G@      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �;@<ݚ)�?             B@        ������������������������       �                     @        �                         �B@�n`���?             ?@       �                       ��yC@      �?
             0@        �                          �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@                                 �?�q�q�?	             .@                               �E@X�Cc�?             ,@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        	                         �?�<ݚ�?             ;@        
                         �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                �7@�q�q�?             8@                                �?�r����?             .@        ������������������������       �                     �?                                 �?؇���X�?
             ,@        ������������������������       �                     @                                 �?"pc�
�?             &@                                  @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                  @r�q��?             @        ������������������������       �                     @                              ��T?@�q�q�?             @        ������������������������       �                     �?                              pf�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  @�q�q�?             "@        ������������������������       �                      @                               �T�E@և���X�?             @        ������������������������       �                     �?        !      "                   ;@      �?             @        ������������������������       �                      @        #      $                �|�>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0M%KK��h2h3h4hVh<�h=Kub������������H�1�N�?oݟ�Kb�?ަ���m�?I�Iψd�?�d�*al�?�YP�9��?9/���?և���X�?�$I�$I�?۶m۶m�?      �?                      �?              �?]t�E�?/�袋.�?      �?      �?      �?                      �?�}A_Ч?�/����?h/�����?�Kh/��?              �?�A�A�?|�W|�W�?333333�?333333�?�q�q�?�q�q�?�?�?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?      �?                      �?�?�������?              �?      �?                      �?/�袋.�?颋.���?�0�0�?��y��y�?v�)�Y7�?#�u�)��?�{a���?������?              �?�������?�������?      �?        �q�q�?�q�q�?              �?�������?�������?      �?                      �?      �?      �?              �?      �?        br1���?�F}g���?KԮD�J�?ە�]���?�������?�������?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?      �?�$I�$I�?�m۶m��?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        �������?�������?              �?      �?        333333�?�������?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        �������?333333�?              �?      �?        �������?ZZZZZZ�?�������?�������?�q�q�?�q�q�?              �?�������?�������?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?ى�؉��?�؉�؉�?      �?      �?              �?      �?        ��.���?t�E]t�?      �?      �?�q�q�?�q�q�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?              �?        |a���?�{a��?/"�Ed�?7����ݼ?�$I�$I�?۶m۶m�?              �?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?��� �l�?=Ѩ�W��?     @�?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�rO#,��?�i��F�?Ṷ�H��?\����չ?�5��P�?(�����?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �q�q�?�q�q�?\���(\�?{�G�z�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?              �?��o��o�?�A�A�?a����?�{a���?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?      �?      �?              �?              �?        333333�?�������?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �1�1�?����?�������?�?n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?              �?        _����z�?
�B�P(�?F]t�E�?F]t�E�?      �?                      �?�������?rY1P»?UUUUUU�?UUUUUU�?              �?      �?      �?۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?              �?      �?      �?      �?        _�^��?z�z��?_�_��?�A�A�?�?�?      �?      �?      �?        ]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?              �?        �������?�?      �?        q=
ףp�?{�G�z�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �|>����?��`0�?���(\��?�z�G��?Q^Cy��?^Cy�5�?F]t�E�?]t�E]�?�q�q�?r�q��?      �?                      �?              �?/�����?B{	�%��?�������?�������?      �?      �?۶m۶m�?�$I�$I�?/�袋.�?F]t�E�?              �?�������?�������?�������?�������?              �?      �?              �?              �?                      �?              �?      �?        �B!��?��{���?      �?      �?�������?UUUUUU�?�������?�������?�$I�$I�?۶m۶m�?              �?;�;��?;�;��?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?��8��8�?�8��8��?              �?�9�s��?�c�1��?      �?      �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?%I�$I��?�m۶m��?              �?      �?              �?              �?        9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?�������?�?      �?        ۶m۶m�?�$I�$I�?      �?        /�袋.�?F]t�E�?�������?�������?              �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?      �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��nhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       f                    �?�,�٧��?�           8�@               M                    �? ْs�?�            pp@              2                   �<@��Y�"��?�            �i@               #                   �8@V�a�� �?6            �U@                                  �?v���a�?+            @R@                                  �2@��<b���?             7@                               P��+@X�Cc�?             ,@        ������������������������       �                     @        	       
                    @      �?             $@        ������������������������       �                     @                                  �-@����X�?             @        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@                                    @H%u��?             I@        ������������������������       �                     4@               "                 ��Y1@z�G�z�?             >@              !                    �?�����H�?             ;@                                  �7@      �?             8@                                  �?���}<S�?             7@        ������������������������       �                     @                                  �5@�t����?             1@        ������������������������       �                      @                                  �6@�<ݚ�?             "@                                �̜!@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?                                @3�@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        $       '                   �9@      �?             ,@        %       &                 hf�2@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        (       -                     @���Q��?             $@        )       ,                   �;@      �?             @        *       +                   �/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        .       1                   �;@      �?             @       /       0                 @3�,@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        3       B                   �B@؞�z�̼?K            @]@       4       7                 ���@ ��WV�?2            �S@        5       6                 �Y�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        8       =                    �?P�Lt�<�?0             S@       9       <                 ��� @@	tbA@�?*            @Q@        :       ;                    �?@4և���?
             ,@       ������������������������       �        	             *@        ������������������������       �                     �?        ������������������������       �                     �K@        >       ?                     @؇���X�?             @        ������������������������       �                     @        @       A                 ���7@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        C       L                     @��-�=��?            �C@       D       E                   @C@@-�_ .�?            �B@        ������������������������       �                     �?        F       K                 �DD@������?             B@        G       J                     �?��S�ۿ?             .@        H       I                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@        ������������������������       �                      @        N       Y                 03�=@�ݜ����?$            �M@        O       T                 �|Y=@�q�q�?             8@       P       S                    +@�t����?             1@        Q       R                    !@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        U       X                 ���8@և���X�?             @       V       W                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        Z       _                     @��R[s�?            �A@        [       ^                     �?      �?              @       \       ]                    $@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        `       a                 X��@@�>����?             ;@       ������������������������       �        	             4@        b       e                 ��p@@����X�?             @        c       d                 ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        g       �                     �?�X�C�?"            |@        h       o                    <@�~�����??            �X@        i       l                    �?�q�q�?             (@        j       k                   �5@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        m       n                  "&d@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        p       �                    �?JyK���?7            �U@       q       r                 ��<:@�M;q��?1            �R@        ������������������������       �                     ,@        s       �                  �>@�-ῃ�?*            �N@        t       w                    �?���|���?             6@        u       v                 ���<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        x       y                 �|Y=@�����?             3@        ������������������������       �                      @        z       �                   @=@������?             1@       {       �                   �J@���|���?             &@       |                        `f�;@�<ݚ�?             "@       }       ~                 �|�?@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �E@x�����?            �C@       �       �                    �?8����?             7@        �       �                 p�w@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                  x#J@�E��ӭ�?             2@       ������������������������       �                     &@        �       �                 `f�N@����X�?             @        ������������������������       �                     @        �       �                 03�S@�q�q�?             @        ������������������������       �                     �?        �       �                 X��@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             0@        ������������������������       �                     @        �       �                 ��#[@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                    �?�8��8��?             (@       �       �                    �?�����H�?             "@       �       �                   @B@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �? ʊ����?�            �u@       �       �                    �?���F6��?�            �r@        �       �                   @@z�G�z�?             9@        �       �                 ���@X�<ݚ�?             "@        �       �                    :@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �5@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     @      �?
             0@        ������������������������       �                     $@        �       �                 �|�;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@�IєX�?�             q@        �       �                    �? ������?R            �_@        ������������������������       �                     6@        �       �                   �7@ pƵHP�?C             Z@        ������������������������       �                    �@@        �       �                   �8@�J�T�?-            �Q@        �       �                 `fF@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��L@����e��?*            �P@       ������������������������       �                    �@@        �       �                    ?@Pa�	�?            �@@       ������������������������       �                     <@        �       �                   �@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @E@����1�?^            @b@       �       �                    �?Xny��?P            �^@        ������������������������       �                     @        �       �                 @3�@�^����?M            �]@        �       �                   �4@      �?              @        ������������������������       �                     �?        �       �                   �A@����X�?             @       ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                 ���"@ףp=
�?G            �[@        �       �                   �2@P�Lt�<�?             C@        �       �                 ��Y @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �@@        �       �                     @4?,R��?/             R@       �       �                   �3@�C��2(�?             F@       �       �                   �C@�t����?             A@       �       �                    &@(;L]n�?             >@        �       �                    5@$�q-�?             *@        ������������������������       ��q�q�?             @        ������������������������       �                     $@        ������������������������       �        
             1@        ������������������������       �      �?             @        ������������������������       �                     $@        �       �                 `�X#@d}h���?             <@        �       �                   �8@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �T)D@���}<S�?             7@       ������������������������       �                     3@        �       �                    ;@      �?             @        ������������������������       �                     �?        �       �                    >@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     8@        �       �                   �C@�n_Y�K�?#             J@       �       �                    �?v ��?            �E@        �       �                 �|Y>@"pc�
�?             &@       �       �                 ��}@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        �       �                 `ff/@     ��?             @@        �       �                     @�C��2(�?             &@        ������������������������       �                      @        �       �                   �*@�����H�?             "@        �       �                    (@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    +@�G��l��?             5@       �       �                    �?����X�?
             ,@        ������������������������       �                     @        �       �                    @�C��2(�?             &@        �       �                     @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������&��jq�?:�g *�?^��{7A�?�U!�/�?______�?�?a���{�?��{a�?�4iҤI�?ٲe˖-�?��Moz��?��,d!�?�m۶m��?%I�$I��?              �?      �?      �?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?���Q��?)\���(�?              �?�������?�������?�q�q�?�q�q�?      �?      �?d!Y�B�?ӛ���7�?              �?�?<<<<<<�?              �?�q�q�?9��8���?�������?�������?              �?      �?              �?      �?              �?      �?              �?                      �?      �?              �?      �?      �?      �?      �?                      �?�������?333333�?      �?      �?      �?      �?              �?      �?                      �?      �?      �?�������?333333�?              �?      �?              �?        �ꡮ?^�^��?;�;��?O��N���?      �?      �?              �?      �?        (�����?���k(�?ہ�v`��?�%~F��?�$I�$I�?n۶m۶�?              �?      �?                      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?        �A�A�?}˷|˷�?к����?S�n0E�?      �?        �q�q�?�q�q�?�?�������?�q�q�?�q�q�?      �?                      �?              �?              �?      �?        �}ylE��?W'u_�?�������?UUUUUU�?�?<<<<<<�?�������?333333�?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?X|�W|��?PuPu�?      �?      �?UUUUUU�?�������?      �?                      �?              �?�Kh/��?h/�����?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �m۶m��?%I�$I��?P�W
���?`)P�W
�?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?333333�?�������?              �?      �?        Ȥx�L��?p��f��?�6�i��?ƒ_,���?      �?        �).�u�?�����?F]t�E�?]t�E]�?UUUUUU�?UUUUUU�?      �?                      �?^Cy�5�?Q^Cy��?      �?        �?xxxxxx�?F]t�E�?]t�E]�?�q�q�?9��8���?      �?      �?      �?                      �?      �?              �?                      �?��o��o�?�A�A�?d!Y�B�?8��Moz�?333333�?�������?      �?                      �?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?۶m۶m�?�$I�$I�?              �?      �?              �?              �?        H6.��=�?�M�V�?�v�ļ�?ogH���?�������?�������?r�q��?�q�q�?      �?      �?              �?      �?        333333�?�������?              �?      �?              �?      �?      �?        �������?UUUUUU�?              �?      �?        �?�?��}��}�?AA�?      �?        'vb'vb�?;�;��?      �?        (�K=�?��V؜?�������?�������?              �?      �?        �>����?|���?      �?        |���?|���?      �?        �������?�������?              �?      �?        �Ν;w��?Ĉ#F��?C��6�S�?�}�K�`�?      �?        u_[4�?W'u_�?      �?      �?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?�������?�������?���k(�?(�����?�������?�������?              �?      �?              �?        �8��8��?r�q��?]t�E�?F]t�E�?<<<<<<�?�?�������?�?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?              �?              �?      �?      �?        I�$I�$�?۶m۶m�?�������?�������?      �?                      �?ӛ���7�?d!Y�B�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ;�;��?ى�؉��?G�w��?qG�w��?F]t�E�?/�袋.�?�������?�������?      �?                      �?      �?              �?      �?]t�E�?F]t�E�?      �?        �q�q�?�q�q�?      �?      �?              �?      �?              �?        1�0��?��y��y�?�$I�$I�?�m۶m��?      �?        F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJXk�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       V                    �?�,�٧��?�           8�@               S                    @��}� �?�            �o@              <                 �|�=@2C�AK0�?�            @n@                                   @*jF���?g            `d@                                    �?0z�(>��?,            �Q@        ������������������������       �                    �A@                                   6@�8��8��?             B@               	                    �?�θ�?	             *@        ������������������������       �                     @        
                           5@�z�G��?             $@        ������������������������       �                     @                                  �;@      �?             @                                 �9@      �?             @                                 �+@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@                                   @(옄��?;             W@                                0CD9@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @               5                    �?      �?4             T@              (                  ��@�2�o�U�?%            �K@                                  �?؇���X�?             <@                                  �?      �?             0@        ������������������������       �                      @                                ���@@4և���?
             ,@        ������������������������       �                     �?        ������������������������       �        	             *@                !                  s@      �?	             (@        ������������������������       �                     @        "       '                    8@�q�q�?             "@       #       $                 ���@؇���X�?             @        ������������������������       �                     @        %       &                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        )       4                 �|�;@|��?���?             ;@       *       3                    3@��Q��?             4@        +       0                    �?�<ݚ�?             "@       ,       -                 �&�)@؇���X�?             @        ������������������������       �                     @        .       /                   �-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        1       2                 �y�+@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        6       ;                 @3�2@HP�s��?             9@        7       8                    �?����X�?             @       ������������������������       �                     @        9       :                   �:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             2@        =       N                   �3@���!���?2            �S@        >       E                   �B@�ՙ/�?             5@       ?       @                     @�8��8��?
             (@       ������������������������       �                     "@        A       B                   �>@�q�q�?             @        ������������������������       �                     �?        C       D                 ��*@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        F       M                 pF4.@�<ݚ�?             "@       G       L                     @      �?              @       H       I                    F@      �?             @        ������������������������       �                      @        J       K                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        O       R                 03�=@ _�@�Y�?"             M@        P       Q                    �?�8��8��?	             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     G@        T       U                    �?r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        W       �                     �?pґ���?!           �|@        X       g                    �?؁sF���?9             Y@        Y       f                 �\@      �?             F@       Z       e                   �H@��Zy�?            �C@       [       d                   @C@������?             >@       \       c                 0��G@D�n�3�?	             3@       ]       `                 X�,@@�q�q�?             (@       ^       _                 �|�;@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        a       b                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     "@        ������������������������       �                     @        h       i                    �?������?%             L@        ������������������������       �                     �?        j       �                 03�U@�b��[��?$            �K@       k       �                   �>@�	j*D�?#             J@       l       w                   �B@�P�*�?             ?@       m       n                 ��I/@D�n�3�?
             3@        ������������������������       �                     @        o       r                 �|Y=@������?             .@        p       q                   �<@      �?             @       ������������������������       �                      @        ������������������������       �                      @        s       v                 `fF<@"pc�
�?             &@       t       u                 �|�?@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        x                           R@r�q��?	             (@       y       z                 `fF:@�C��2(�?             &@        ������������������������       �                     @        {       ~                 `f�;@      �?              @       |       }                   @I@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���L@؇���X�?             5@       �       �                 `fFJ@z�G�z�?             .@       �       �                   �A@�C��2(�?	             &@        ������������������������       �                     @        �       �                 ��yC@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    7@      �?             @        ������������������������       �                     �?        �       �                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?0y����?�            Pv@       �       �                 0C�E@؅�q(�?�            �r@       �       �                    ,@@�z���?�            �r@        �       �                    '@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �E@�U�:��?�            pr@       �       �                 ���@�?�(|�?�            pp@        ������������������������       �                     ;@        �       �                     @����>�?�            �m@        �       �                   �C@4��?�?             J@       �       �                    5@ �q�q�?             H@        �       �                   �'@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                 �|�=@ qP��B�?            �E@       �       �                    �?P���Q�?             4@        ������������������������       �                     @        �       �                 �|Y=@�IєX�?             1@       ������������������������       �        
             0@        ������������������������       �                     �?        ������������������������       �                     7@        �       �                    4@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q��/��?|             g@        �       �                   �+@      �?             @@       �       �                   �6@ףp=
�?             >@        ������������������������       �                      @        �       �                 ���@h�����?             <@        ������������������������       �                     $@        �       �                 �|Y?@�X�<ݺ?	             2@       �       �                   @@@4և���?             ,@       �       �                 �|=@      �?              @        ������������������������       �                     @        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���@�KM�]�?j             c@        ������������������������       �                      @        �       �                   @C@���Lͩ�?i            �b@       �       �                 �|�=@T�n��?e             b@       �       �                 м�5@�&/�E�?V             _@       �       �                 @3�!@�.ߴ#�?T            �^@       �       �                    �?8v�YeK�?D            �W@        �       �                  ��@      �?
             0@        ������������������������       �                     @        �       �                 ��(@ףp=
�?             $@       �       �                 �|Y=@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �0@86��Z�?:            �S@        ������������������������       ��q�q�?             @        �       �                   �:@�}�+r��?8             S@       �       �                 @3�@����?�?!            �F@       ������������������������       �                     >@        �       �                 0S5 @��S�ۿ?             .@       �       �                   �4@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �;@��a�n`�?             ?@        �       �                 �� @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �&B@@4և���?             <@        �       �                 ��,@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|Y=@`2U0*��?             9@        ������������������������       �                     @        �       �                 ��) @���7�?             6@       ������������������������       �                     3@        �       �                 pf� @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ;@        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �?@z�G�z�?             4@        �       �                 �?�@և���X�?             @        ������������������������       �                     @        �       �                 @3�@      �?             @        ������������������������       �                      @        �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @@@$�q-�?
             *@       �       �                 ��I @      �?              @       �       �                 �?�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    D@      �?             @       �       �                 ��	0@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @@        �       �                 ��?P@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �                          @����0�?&             K@        �       �                     @     ��?             0@       ������������������������       �                     "@        �                          @և���X�?             @       �                        8#8@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                              �|Y>@�S����?             C@                             �̌4@�θ�?             :@                              ��\"@      �?              @        ������������������������       �                     �?                              032@؇���X�?             @       ������������������������       �                     @        	      
                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �        	             (@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������&��jq�?:�g *�?�@ �?��~����?3(&ޏ�?�zv��?��0��?~��g*�?H���@��?�ԓ�ۥ�?              �?UUUUUU�?UUUUUU�?�؉�؉�?ى�؉��?              �?333333�?ffffff�?              �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?ӛ���7�?���,d�?UUUUUU�?�������?              �?      �?              �?      �?�S�<%��?־a��?�$I�$I�?۶m۶m�?      �?      �?              �?�$I�$I�?n۶m۶�?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?        	�%����?{	�%���?�������?ffffff�?�q�q�?9��8���?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?              �?                      �?q=
ףp�?{�G�z�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        T:�g *�?��	�Z�?�a�a�?�<��<��?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        9��8���?�q�q�?      �?      �?      �?      �?      �?              �?      �?              �?      �?              �?                      �?�{a���?#,�4�r�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?UUUUUU�?              �?      �?        �����?J�!����?�z�G��?=
ףp=�?      �?      �?\��[���?� � �?�?wwwwww�?(������?l(�����?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?        �������?333333�?              �?      �?                      �?              �?      �?              �?        I�$I�$�?n۶m۶�?      �?        � O	��?־a��?vb'vb'�?;�;��?�RJ)���?�Zk����?(������?l(�����?      �?        �?wwwwww�?      �?      �?              �?      �?        F]t�E�?/�袋.�?�������?333333�?      �?                      �?              �?�������?UUUUUU�?]t�E�?F]t�E�?      �?              �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?                      �?۶m۶m�?�$I�$I�?�������?�������?]t�E�?F]t�E�?      �?        �������?UUUUUU�?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?�5�5�?gZ{���?e�,%l��?��y���?}0T�1�?UUUUUU�?UUUUUU�?      �?                      �?�A�I�?�pR�屵?��X�J��?]`;e�U�?      �?        _[4��?'u_�?�N��N��?ى�؉��?�������?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?        ��}A�?�}A_З?ffffff�?�������?      �?        �?�?      �?                      �?      �?              �?      �?              �?      �?        �B����?��Mozӻ?      �?      �?�������?�������?              �?�m۶m��?�$I�$I�?      �?        ��8��8�?�q�q�?n۶m۶�?�$I�$I�?      �?      �?      �?        �������?�������?      �?              �?              �?      �?              �?      �?        �k(���?(�����?              �?�6�i�?�K~��?�8��8��?�8��8��?2�c�1�?�s�9�?�K�`m�?XG��).�?��sK���?�a�+�?      �?      �?      �?        �������?�������?�q�q�?�q�q�?              �?      �?              �?        �Z܄��?h *�3�?UUUUUU�?UUUUUU�?�5��P�?(�����?��I��I�?l�l��?      �?        �������?�?      �?      �?              �?      �?              �?        �s�9��?�c�1Ƹ?UUUUUU�?UUUUUU�?      �?                      �?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?���Q��?{�G�z�?      �?        �.�袋�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?        �������?�������?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?      �?      �?                      �?�؉�؉�?;�;��?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?              �?      �?�������?333333�?      �?      �?      �?              �?              �?        333333�?�������?              �?      �?        �Kh/���?Lh/����?      �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?                      �?(������?^Cy�5�?ى�؉��?�؉�؉�?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ0��JhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                  x#J@ʻ�J��?�           8�@              I                     @��+7��?y           ��@                                   @�1�x��?�            �j@        ������������������������       �                      @               6                    �?��+1�+�?�            �i@              3                  �>@�����C�?d             d@                                  �?�7�֥��?R            @`@                                    �?(L���?            �E@        	       
                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                  �I@$G$n��?            �B@                                 �;@�����H�?             B@                                   9@      �?             (@       ������������������������       �                     @                                ��m1@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @                                  �B@ �q�q�?             8@       ������������������������       �        	             1@                                  �C@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               (                     �?�=C|F�?:            �U@                                  �<@�q�q�?             8@        ������������������������       �                      @               !                    �?���!pc�?             6@                                �|�=@      �?             @        ������������������������       �                      @                                 `f&;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        "       '                    R@r�q��?             2@       #       $                   �G@�t����?
             1@        ������������������������       �                     "@        %       &                   @L@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        )       ,                    4@���N8�?*            �O@        *       +                   �2@�<ݚ�?             "@        ������������������������       �                     @        ������������������������       ��q�q�?             @        -       2                 �|�=@@3����?&             K@        .       /                    �?���N8�?             5@        ������������������������       �                     @        0       1                 �|Y=@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                    �@@        4       5                    �?�חF�P�?             ?@        ������������������������       �                     @        ������������������������       �                     :@        7       H                 �%D@      �?             F@       8       9                     �?>��C��?            �E@        ������������������������       �                     �?        :       ;                    �?d}h���?             E@        ������������������������       �                     �?        <       E                   �:@� ��1�?            �D@       =       D                    @�X����?             6@       >       ?                    �?��Q��?             4@       ������������������������       �        
             &@        @       C                    �?�<ݚ�?             "@       A       B                    1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        F       G                   �A@�}�+r��?
             3@       ������������������������       �        	             2@        ������������������������       �                     �?        ������������������������       �                     �?        J       �                    �?"pc�
�?�            x@        K       �                 �|�=@����3��?D             Z@       L       �                   0:@��C���?<            �W@       M       b                    �?�L��7Q�?9            @V@        N       ]                    �?     ��?             @@        O       \                 `�@1@�eP*L��?	             &@       P       Q                   �"@      �?              @        ������������������������       �                     �?        R       Y                    �?����X�?             @       S       X                    �?z�G�z�?             @       T       U                 �|6@      �?             @        ������������������������       �                     �?        V       W                 ��%@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        Z       [                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ^       _                 ���@�����?             5@        ������������������������       �                     �?        `       a                    �?P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        c       x                    �?�MWl��?#            �L@        d       o                   �<@���Q��?             9@       e       l                 �0@����X�?	             ,@       f       g                ��k$@"pc�
�?             &@        ������������������������       �                     �?        h       k                 ���@ףp=
�?             $@        i       j                 ��y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        m       n                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        p       w                    �?�eP*L��?             &@       q       r                 �|Y=@      �?              @        ������������������������       �                     �?        s       t                 ���@����X�?             @        ������������������������       �                     �?        u       v                   @@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     @        y       |                 �|Y=@     ��?             @@        z       {                    ;@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        }       �                   `3@@4և���?             <@       ~                        ���@ 7���B�?             ;@        ������������������������       �                     @        �       �                 ��(@�nkK�?             7@       ������������������������       ��}�+r��?
             3@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    @�n3�F��?�            �q@        �       �                 @3�4@���|���?
             &@        ������������������������       �                      @        �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                 `f�:@�q�q�?             @        ������������������������       �                     �?        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �̌4@�Aʑ���?�            �p@       �       �                 03c4@<���D�?�            �l@       �       �                    �?��O���?�            �l@        �       �                    �?X�<ݚ�?             B@       �       �                 pf�@և���X�?            �A@        ������������������������       �                     @        �       �                 @3�@�q�q�?             >@        �       �                    6@և���X�?             @        ������������������������       �                      @        �       �                   �9@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y=@��+7��?             7@        �       �                  �M$@�8��8��?             (@        �       �                    3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��� @�eP*L��?             &@        ������������������������       �                      @        �       �                   �>@X�<ݚ�?             "@        ������������������������       �                     @        �       �                  SE"@�q�q�?             @        ������������������������       �                     �?        �       �                   �@@z�G�z�?             @        ������������������������       �                      @        �       �                 `f�/@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�0p<���?s             h@       �       �                   �2@Ȥ4"��?o             g@        ������������������������       �                     3@        �       �                   @4@`�f��?g            �d@        �       �                 0S5 @؇���X�?             5@       �       �                 �?�@      �?             (@        ������������������������       �                     @        �       �                 @3�@և���X�?             @        ������������������������       �                      @        �       �                   �3@z�G�z�?             @       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     "@        �       �                 ��) @ )�y���?X             b@       �       �                 ��@ f^8���?B            �Y@        ������������������������       �                     >@        �       �                    ?@���(-�?/            @R@       �       �                 �?$@�O4R���?#            �J@        ������������������������       ��q�q�?             @        ������������������������       �        !             I@        �       �                 @3�@ףp=
�?             4@       �       �                 �&B@8�Z$���?             *@        ������������������������       �                     @        �       �                   �A@����X�?             @       �       �                   �@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                    ?@���H��?             E@       �       �                 �|�=@�חF�P�?             ?@       �       �                 pf� @ܷ��?��?             =@        ������������������������       �                     @        ������������������������       �                     :@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @        �       �                    5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �C@        �                          O@
�ۓQ{�?J            @\@       �       �                    �?����|e�?G             [@       �       �                     @�.ߴ#�?,            �N@       ������������������������       �        *             M@        ������������������������       �                     @        �       �                 `�>P@z�J��?            �G@        �       �                      @"pc�
�?             &@       �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �                    7@      �?             @        ������������������������       �                     �?        �       �                 `f�K@�q�q�?             @       �       �                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?             B@       �       �                 p�w@և���X�?
             5@       �       �                  �}S@      �?             2@        ������������������������       �                      @        �       �                    �?     ��?             0@       �       �                    �?�	j*D�?             *@       �       �                   �8@�q�q�?             (@        ������������������������       �                     @        �       �                 �|Y;@z�G�z�?             @        ������������������������       �                      @        �       �                 0�c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �                          �?z�G�z�?	             .@       �                           �?$�q-�?             *@       �       �                 X��@@ףp=
�?             $@        ������������������������       �                     @        �       �                 03�U@r�q��?             @        ������������������������       �                     @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������"N���I�?�c�~`l�?zӛ����?Y�B��?8��n�?���"��?      �?        ��5)[��?ٚ��I��?��J1Aw�?��j�}�?�B/�B/�?z�z��?w�qG��?⎸#��?UUUUUU�?�������?      �?                      �?���L�?к����?�q�q�?�q�q�?      �?      �?              �?۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?�������?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?        �C��:��?J��/�?UUUUUU�?UUUUUU�?              �?F]t�E�?t�E]t�?      �?      �?              �?      �?      �?              �?      �?        �������?UUUUUU�?<<<<<<�?�?      �?              �?      �?              �?      �?                      �?��y��y�?�a�a�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?���Kh�?h/�����?��y��y�?�a�a�?      �?        �������?�?      �?                      �?      �?        �Zk����?��RJ)��?              �?      �?              �?      �?qG�w��?$�;��?      �?        ۶m۶m�?I�$I�$�?      �?        ������?������?]t�E]�?�E]t��?ffffff�?�������?              �?9��8���?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?(�����?�5��P�?              �?      �?              �?        /�袋.�?F]t�E�?��N��N�?'vb'vb�?L� &W�?g���Q��?%+Y�JV�?��MmjS�?      �?      �?]t�E�?t�E]t�?      �?      �?              �?�m۶m��?�$I�$I�?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?                      �?�a�a�?=��<���?      �?        �������?ffffff�?              �?      �?        :��,���?�YLg1�?333333�?�������?�m۶m��?�$I�$I�?/�袋.�?F]t�E�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?]t�E�?t�E]t�?      �?      �?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?                      �?      �?      �?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?	�%����?h/�����?      �?        �Mozӛ�?d!Y�B�?�5��P�?(�����?      �?                      �?      �?              �?        �t�k[�?[��,'�?]t�E]�?F]t�E�?              �?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        ���u��?Ũ�oS��?|���?|���?���!:�?D����.�?r�q��?�q�q�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?                      �?zӛ����?Y�B��?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?        t�E]t�?]t�E�?      �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?��3-�?�O�l.�?���y��?�cxq�?      �?        ��(��?�7�:���?۶m۶m�?�$I�$I�?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?      �?      �?      �?              �?        q��<�?����?�?H%�e�?��VCӝ?      �?        ��իW��?�P�B�
�?:�&oe�?�x+�R�?UUUUUU�?UUUUUU�?      �?        �������?�������?;�;��?;�;��?      �?        �m۶m��?�$I�$I�?�������?�������?              �?      �?              �?      �?      �?        �0�0�?��y��y�?�Zk����?��RJ)��?��=���?a���{�?              �?      �?                      �?      �?              �?              �?      �?              �?      �?              �?        ��Ź��?2�s�8�?	�%����?����K�?XG��).�?�K�`m�?              �?      �?        }g���Q�?AL� &W�?F]t�E�?/�袋.�?�q�q�?9��8���?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?�������?�������?۶m۶m�?�$I�$I�?      �?      �?              �?      �?      �?vb'vb'�?;�;��?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?�������?�������?�؉�؉�?;�;��?�������?�������?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJڡWhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       L                 @3�"@�����?�           8�@                                   �?H�g�}N�?�            q@                                   �?�	j*D�?             :@                                 �6@�q�q�?             8@        ������������������������       �                     &@                                �?�@�n_Y�K�?	             *@              
                    �?�<ݚ�?             "@               	                 �&�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                  �8@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                               ��k @@�?��K�?�            �n@        ������������������������       �                     �?                                ���@,��w�?�            �n@        ������������������������       �                    �G@               K                   �C@�`��H �?z            �h@                               ��@��F��9�?n             f@        ������������������������       �                      @               "                 �Y�@�#-���?m            �e@                                ���@�d�����?             3@                                �|�9@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                                  �5@���Q��?             $@        ������������������������       �                      @                                �|�:@      �?              @        ������������������������       �                      @                !                 �|�=@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        #       2                 �?�@ ��Ou��?b            �c@       $       %                   �<@�==Q�P�?;            �W@        ������������������������       �                    �G@        &       1                 �Yu@      �?             H@       '       0                 ��]@ףp=
�?             >@       (       )                 ���@ 	��p�?             =@        ������������������������       �                     &@        *       +                 �|Y=@�����H�?             2@        ������������������������       �                     �?        ,       -                    �?�IєX�?
             1@       ������������������������       �                     *@        .       /                 �|Y?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             2@        3       4                    �?Xny��?'            �N@        ������������������������       �                      @        5       D                 0SE @�^����?&            �M@       6       C                 ��) @8�Z$���?            �C@       7       :                   �3@������?            �B@        8       9                   �1@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ;       B                   �B@      �?             @@       <       A                 @3�@(;L]n�?             >@        =       >                   �=@      �?              @        ������������������������       �                     @        ?       @                   �?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     6@        ������������������������       �      �?              @        ������������������������       �                      @        E       F                 @Q!@P���Q�?             4@        ������������������������       �                      @        G       J                 @3�!@�8��8��?             (@       H       I                   �:@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     6@        M       �                    �?ȱma���?           `{@        N       y                    �?v���6h�?�            `j@       O       h                     @�����8�?H            @]@       P       g                 03�>@,���$�?;            @X@       Q       X                   �B@L紂P�?            �I@       R       W                   �9@      �?             @@        S       T                   �7@z�G�z�?             @       ������������������������       �                     @        U       V                   �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ;@        Y       \                     �?�����?             3@        Z       [                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ]       f                    L@�n_Y�K�?             *@       ^       c                    5@���!pc�?             &@       _       b                   �*@؇���X�?             @        `       a                   �'@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        d       e                   �E@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     G@        i       x                 ���1@�G�z��?             4@       j       k                   �#@     ��?             0@        ������������������������       �                     @        l       m                   @0@�n_Y�K�?
             *@        ������������������������       �                      @        n       o                    �?���!pc�?	             &@        ������������������������       �                     �?        p       q                    �?z�G�z�?             $@        ������������������������       �                     �?        r       s                 Ь�#@�<ݚ�?             "@        ������������������������       �                     �?        t       w                 ��&@      �?              @        u       v                 �[$@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        z                            @�7����?9            �W@       {       |                 ���a@@3����?              K@       ������������������������       �                     E@        }       ~                    '@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?      �?             D@        �       �                 `�@1@���Q��?             $@       �       �                    �?؇���X�?             @       �       �                 P��+@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @d��0u��?             >@        �       �                    �?؇���X�?             @       �       �                     @r�q��?             @        ������������������������       �                     @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�2@��<b���?             7@        �       �                    :@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @�X�<ݺ?             2@       ������������������������       �        	             .@        �       �                 ���A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @(����?�            `l@        �       �                 �Q��?p�ݯ��?             3@        ������������������������       �                     @        �       �                   �;@��S���?             .@        ������������������������       �                     @        �       �                    @���|���?             &@        �       �                 �D,C@r�q��?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                      @���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                 ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�θ�?�             j@       �       �                     �?����|e�?n            @d@        �       �                   �;@:%�[��?2            �Q@        �       �                   �8@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                  x#J@f���M�?+             O@       �       �                  �>@���3�E�?#             J@       �       �                    �?l��[B��?             =@        �       �                   @G@���Q��?             $@       �       �                   @@@      �?              @       �       �                 �|�=@�q�q�?             @       �       �                 �ܵ<@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 �|Y=@�\��N��?             3@        ������������������������       �                      @        �       �                   @=@j���� �?             1@       �       �                 ��$:@�z�G��?             $@        ������������������������       �                     @        �       �                    D@      �?             @        ������������������������       �                     �?        �       �                 `f�;@���Q��?             @       �       �                   @G@      �?             @        ������������������������       �                     �?        �       �                   @L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �B@�nkK�?             7@        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                 �TaA@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                 �|Y>@�z�G��?             $@        ������������������������       �                      @        �       �                    �?      �?              @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @Ĝ�oV4�?<            �V@       �       �                   �@@�}�+r��?%            �L@       �       �                    &@�?�|�?            �B@        �       �                   �5@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     ?@        �       �                   �A@ףp=
�?             4@        �       �                    1@����X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �        	             *@        �       �                    9@������?             A@        �       �                    ,@$�q-�?	             *@        �       �                 �y.@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 �T)D@�q�q�?             5@       �       �                 pF�'@�d�����?             3@        �       �                   �?@      �?             @       �       �                   �<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   @;@8�Z$���?             *@        �       �                 �0@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        �       �                     �?�3Ea�$�?             G@        �       �                   �7@      �?	             0@        ������������������������       �                     @        ������������������������       �                     (@        �                           �?r�q��?             >@        �       �                     @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                 #@HP�s��?             9@                                 �?�q�q�?             @        ������������������������       �                     @                                  @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�����������������?��܍��?|��{���?���?;�;��?vb'vb'�?UUUUUU�?UUUUUU�?              �?;�;��?ى�؉��?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?              �?�����?~*! 秲?              �?�-�����?��鰱?      �?        R@�O.D�?m�큍޵?k��2��?�L;k��?              �?�A�A�?_�_�?Cy�5��?y�5���?�q�q�?�q�q�?              �?      �?        333333�?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?        .��-���?�i�i�?��%N��?�a�+�?      �?              �?      �?�������?�������?������?�{a���?      �?        �q�q�?�q�q�?              �?�?�?      �?              �?      �?              �?      �?                      �?      �?        C��6�S�?�}�K�`�?      �?        u_[4�?W'u_�?;�;��?;�;��?��g�`��?к����?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?�������?�?      �?      �?      �?              �?      �?              �?      �?              �?              �?      �?              �?ffffff�?�������?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?      �?              �?        ��{���?��.��?�iP�z�?�%�k]��?���?�������?���fy�?�,O"Ӱ�?�������?�������?      �?      �?�������?�������?              �?      �?      �?      �?                      �?              �?^Cy�5�?Q^Cy��?UUUUUU�?�������?      �?                      �?ى�؉��?;�;��?t�E]t�?F]t�E�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?              �?                      �?�������?�������?      �?      �?              �?ى�؉��?;�;��?      �?        t�E]t�?F]t�E�?      �?        �������?�������?              �?�q�q�?9��8���?      �?              �?      �?      �?      �?              �?      �?                      �?      �?        G}g����?]AL� &�?h/�����?���Kh�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?333333�?�������?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?                      �?DDDDDD�?wwwwww�?�$I�$I�?۶m۶m�?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?��,d!�?��Moz��?�������?�������?              �?      �?        ��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �]/����?�D�����?Cy�5��?^Cy�5�?              �?�������?�?              �?]t�E]�?F]t�E�?�������?UUUUUU�?      �?      �?              �?      �?              �?        �������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?ى�؉��?�؉�؉�?����K�?	�%����?+l$Za�?�'�K=�?UUUUUU�?UUUUUU�?      �?                      �?��RJ)��?��Zk���?O��N���?b'vb'v�?���=��?GX�i���?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?333333�?�������?      �?                      �?      �?                      �?      �?        �5��P�?y�5���?      �?        ZZZZZZ�?�������?ffffff�?333333�?      �?              �?      �?              �?333333�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�Mozӛ�?d!Y�B�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?        333333�?ffffff�?      �?              �?      �?      �?      �?              �?      �?                      �?�!�!�?����?�5��P�?(�����?*�Y7�"�?к����?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        �������?�������?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?        xxxxxx�?�?�؉�؉�?;�;��?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?Cy�5��?y�5���?      �?      �?      �?      �?      �?                      �?      �?        ;�;��?;�;��?      �?      �?      �?                      �?      �?                      �?����7��?��,d!�?      �?      �?              �?      �?        �������?UUUUUU�?�������?333333�?      �?                      �?q=
ףp�?{�G�z�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:d�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                  x#J@�4�O��?�           8�@              S                    �?
����y�?z           �@                                    @v�X��?r             f@                                   �?�����H�?-             R@        ������������������������       �                     &@                                   L@(��+�?&            �N@                                  �?��ϭ�*�?%             M@                                 �;@д>��C�?             =@        	       
                   �'@և���X�?             @        ������������������������       �                      @                                  �5@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                 ��9@�C��2(�?             6@       ������������������������       �        
             .@                                   D@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     =@        ������������������������       �                     @                                 ��@
j*D>�?E             Z@                                ��@���7�?             6@       ������������������������       �        
             ,@                                   @      �?              @                                  �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               N                    @�W����?5            �T@              M                   @D@�EH,���?0            �R@              0                    �?��z4���?-            @Q@                '                    �?�<ݚ�?             2@        !       &                 pF�-@�C��2(�?             &@        "       #                 �&�)@r�q��?             @        ������������������������       �                      @        $       %                   �-@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        (       )                    @և���X�?             @        ������������������������       �                      @        *       +                    5@���Q��?             @        ������������������������       �                      @        ,       -                 �|�:@�q�q�?             @        ������������������������       �                     �?        .       /                  S�2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       L                 �|�=@��.k���?             �I@       2       A                 ��Y1@�zv�X�?             F@       3       >                    �?      �?             :@       4       9                  �#@D�n�3�?             3@       5       6                   �9@r�q��?             (@       ������������������������       �                     "@        7       8                 �|�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        :       ;                 @3�,@؇���X�?             @        ������������������������       �                     @        <       =                 �|�;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ?       @                    :@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        B       C                 �̌5@�<ݚ�?             2@        ������������������������       �                     @        D       E                    �?�q�q�?	             (@        ������������������������       �                      @        F       K                    @���Q��?             $@        G       H                 `f�:@z�G�z�?             @        ������������������������       �                      @        I       J                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        O       P                    @؇���X�?             @        ������������������������       �                     �?        Q       R                   @C@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        T       �                    �?�/��Y��?           {@       U       p                    �?�@���?�            �w@        V       c                     @�LQ�1	�?!             G@        W       b                     �?������?             1@       X       Y                 �|�;@�q�q�?
             (@        ������������������������       �                     �?        Z       [                 `f&;@���!pc�?	             &@        ������������������������       �                     �?        \       ]                    C@z�G�z�?             $@        ������������������������       �                     @        ^       _                  �>@���Q��?             @        ������������������������       �                      @        `       a                 �D D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        d       o                 �0@�f7�z�?             =@       e       f                   �7@��>4և�?             <@        ������������������������       �                      @        g       h                   �<@R���Q�?             4@        ������������������������       �                     @        i       j                 ���@d}h���?             ,@        ������������������������       �                     @        k       l                 �|Y=@�q�q�?             "@        ������������������������       �                      @        m       n                   @@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        q       �                     �?������?�            �t@        r       s                   �;@>��C��?            �E@        ������������������������       �                     �?        t       �                    R@d}h���?             E@       u       ~                    A@� ��1�?            �D@        v       }                   �>@�KM�]�?             3@        w       |                   @>@�<ݚ�?             "@       x       y                 `f�;@      �?              @        ������������������������       �                     @        z       {                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@               �                   �J@���!pc�?             6@       �       �                 �T!@@      �?
             0@       �       �                   �=@�eP*L��?             &@       �       �                   �9@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                 03k:@      �?              @        ������������������������       �                     �?        �       �                 `f�;@և���X�?             @       �       �                   @G@      �?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @E@�8��8N�?�             r@       �       �                    �?�L���?�            0p@        �       �                 �|Y=@PN��T'�?             ;@        ������������������������       �                     �?        �       �                 X��A@ȵHPS!�?             :@       �       �                   `3@H%u��?             9@       �       �                 ��(@���N8�?             5@       �       �                 ���@$�q-�?	             *@        ������������������������       �                      @        ������������������������       ��C��2(�?             &@        ������������������������       �                      @        �       �                 03�7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �>@Z0Rb�?�             m@       �       �                     @�tVV�?k            �g@        �       �                    &@P�Lt�<�?             C@        �       �                    @�X�<ݺ?
             2@        ������������������������       �                     "@        �       �                    5@�����H�?             "@        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        
             4@        �       �                 �?�@Х-��ٹ?W            �b@       ������������������������       �        ,            �S@        �       �                 @3�@�����H�?+             R@        �       �                   �4@�q�q�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        �       �                 ���#@�[|x��?'            �O@       �       �                   �:@�����H�?            �F@        �       �                   �3@�nkK�?             7@       �       �                   �2@�8��8��?             (@       ������������������������       �                     $@        ������������������������       �      �?              @        ������������������������       �                     &@        �       �                 ��) @"pc�
�?             6@       ������������������������       �        
             .@        �       �                   �;@և���X�?             @        ������������������������       �                     �?        �       �                   �<@      �?             @        ������������������������       �                     �?        �       �                 �|Y=@���Q��?             @        ������������������������       �                     �?        �       �                 pf� @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             2@        �       �                   @@@"pc�
�?             F@        �       �                   �?@      �?              @        �       �                 pff@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 P�@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �?�@�8��8��?             B@        ������������������������       �                     .@        �       �                     @؇���X�?             5@       �       �                   �3@ףp=
�?             $@        �       �                 `fF)@      �?             @        ������������������������       �                     �?        �       �                   @D@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �B@"pc�
�?             &@       ������������������������       �                     @        �       �                   @D@���Q��?             @       �       �                 ��	0@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     =@        �       �                    @������?             L@        �       �                     @���y4F�?             3@        ������������������������       �                     @        �       �                    �?������?	             .@       �       �                    �?�z�G��?             $@        ������������������������       �                     �?        �       �                    �?�q�q�?             "@        ������������������������       �                     �?        �       �                 pf�0@      �?              @        ������������������������       �                     @        ������������������������       �                      @        �       �                    @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?������?            �B@        �       �                     @���Q��?             @        ������������������������       �                     �?        �       �                   �2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    $@      �?             @@        �       �                    �?����X�?             @       �       �                     @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     9@        �       �                    �?t�F�}�?D            �Y@       �       �                    �?l�b�G��?&            �L@       ������������������������       �                    �F@        �       �                    �?�q�q�?             (@        ������������������������       �                     �?        �       �                 �|�:@���|���?             &@        ������������������������       �                     @        �       �                     @և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       
                   <@��S���?            �F@               	                    @������?
             .@                              "�h@�	j*D�?	             *@                                 �?"pc�
�?             &@                              �}S@ףp=
�?             $@       ������������������������       �                     @                              0�HU@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                              X�,@@�q�q�?             >@        ������������������������       �                     @                              �UcV@\X��t�?             7@                                �H@�q�q�?             (@                               �G@�z�G��?             $@                                �E@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                �D@���!pc�?             &@                                 �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                              ��^@      �?              @       ������������������������       �                     @                                �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������X�>�?2�N����?g��4�?3�����?颋.���?�.�袋�?�q�q�?�q�q�?              �?;ڼOq��?q�����?|a���?����=�?|a���?a���{�?۶m۶m�?�$I�$I�?              �?333333�?�������?              �?      �?        F]t�E�?]t�E�?              �?�$I�$I�?�m۶m��?              �?      �?                      �?      �?        ;�;��?b'vb'v�?F]t�E�?�.�袋�?              �?      �?      �?      �?      �?              �?      �?                      �?��|���?p>�cp�?�_,�Œ�?7�i�6�?̵s���?%~F���?�q�q�?9��8���?F]t�E�?]t�E�?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?�?��.���?�袋.��?      �?      �?l(�����?(������?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?�$I�$I�?�m۶m��?              �?      �?        9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?        333333�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?              �?      �?        N<�U�?�����?�ȘW��?�9CE�?Nozӛ��?d!Y�B�?xxxxxx�?�?UUUUUU�?UUUUUU�?              �?F]t�E�?t�E]t�?              �?�������?�������?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        O#,�4��?a���{�?۶m۶m�?I�$I�$�?              �?333333�?333333�?      �?        I�$I�$�?۶m۶m�?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?t�� �?@�_���?$�;��?qG�w��?              �?I�$I�$�?۶m۶m�?������?������?�k(���?(�����?9��8���?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        F]t�E�?t�E]t�?      �?      �?]t�E�?t�E]t�?r�q��?�q�q�?      �?              �?      �?              �?�$I�$I�?۶m۶m�?      �?      �?333333�?�������?              �?      �?                      �?      �?              �?                      �?�������?�������?}���g�?L�Ϻ��?&���^B�?h/�����?              �?��N��N�?�؉�؉�?)\���(�?���Q��?��y��y�?�a�a�?�؉�؉�?;�;��?      �?        ]t�E�?F]t�E�?      �?              �?      �?              �?      �?              �?        �{a���?O#,�4²?ڨ�l�w�?br1���?���k(�?(�����?��8��8�?�q�q�?      �?        �q�q�?�q�q�?      �?      �?      �?              �?        K~��K�?O贁N�?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?      �?      �?        ]�u]�u�?EQEQ�?�q�q�?�q�q�?�Mozӛ�?d!Y�B�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        /�袋.�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?              �?      �?      �?      �?        �������?333333�?              �?      �?      �?              �?      �?              �?        /�袋.�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?              �?      �?        UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        /�袋.�?F]t�E�?      �?        333333�?�������?      �?      �?              �?      �?              �?              �?        I�$I�$�?n۶m۶�?(������?6��P^C�?              �?�?wwwwww�?333333�?ffffff�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?�������?              �?      �?        ��g�`��?к����?333333�?�������?      �?              �?      �?      �?                      �?      �?      �?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?              �?        �������?777777�?p�}��?�Gp��?              �?UUUUUU�?UUUUUU�?              �?F]t�E�?]t�E]�?              �?�$I�$I�?۶m۶m�?              �?      �?        �?�������?�?wwwwww�?;�;��?vb'vb'�?F]t�E�?/�袋.�?�������?�������?              �?      �?      �?      �?                      �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?        !Y�B�?��Moz��?�������?�������?333333�?ffffff�?      �?      �?              �?      �?                      �?      �?        F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?              �?      �?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�I]fhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       z                 ��K.@�L*�<�?�           8�@                                 �,@����?�             x@        ������������������������       �                     @                                03�@.|S͸�?�            �w@        ������������������������       �                    �G@               %                     @<���3��?�            �t@                                   �?�r*e���?,            �R@               	                 `f�)@���}<S�?             7@        ������������������������       �                      @        
                          �*@�r����?
             .@                                  �?"pc�
�?             &@                                  :@�<ݚ�?             "@        ������������������������       �                     �?                                   B@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �?�t����?            �I@        ������������������������       �                     @                                  �(@��E�B��?            �G@        ������������������������       �                     1@               $                   �*@z�G�z�?             >@                                  @@V�a�� �?             =@                               �|�=@��S�ۿ?	             .@                               �|�<@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @               #                   �F@X�Cc�?             ,@              "                   @D@      �?             $@               !                   @B@և���X�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        &       y                   @@@<�I<���?�             p@       '       >                    �?"M�ŋ��?�             k@        (       -                 ��@
j*D>�?!             J@        )       *                 ���@�KM�]�?             3@       ������������������������       �                     &@        +       ,                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        .       /                    �?����e��?            �@@        ������������������������       �                     @        0       =                    �?���>4��?             <@       1       2                    �?���Q��?             9@        ������������������������       �                     @        3       <                 �|�=@�X����?             6@       4       7                    3@���y4F�?             3@        5       6                 ��!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        8       9                   �9@      �?	             0@       ������������������������       �                     (@        :       ;                 @3�@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ?       T                 �?$@<���D�?b            �d@        @       Q                 ��@��.��?&            �N@       A       D                   �7@      �?#             L@        B       C                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        E       F                   �<@ i���t�?            �H@        ������������������������       �                     $@        G       N                  s�@�ݜ�?            �C@       H       M                    �?P���Q�?             4@        I       J                 ���@�����H�?             "@        ������������������������       �                     @        K       L                 �|�=@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     &@        O       P                 �|Y=@���y4F�?
             3@        ������������������������       �                     �?        ������������������������       �r�q��?	             2@        R       S                 �|Y8@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        U       Z                    �?4��?�?<             Z@        V       Y                 ��Y&@�q�q�?             @       W       X                 �|Y=@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        [       ^                   �2@Hm_!'1�?8            �X@        \       ]                   �1@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        _       `                    �?���L��?3            �V@        ������������������������       �                     �?        a       r                 �|�=@��S�ۿ?2            �V@       b       c                 �?�@H�!b	�?+            @T@        ������������������������       �                     =@        d       g                   �4@$�q-�?             J@        e       f                 @3�@8�Z$���?             *@        ������������������������       �      �?             @        ������������������������       �                     "@        h       i                 ��) @�7��?            �C@       ������������������������       �                     =@        j       k                   �<@z�G�z�?             $@        ������������������������       �                     @        l       q                    (@���Q��?             @       m       n                 `��!@�q�q�?             @        ������������������������       �                     �?        o       p                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        s       t                   �@�<ݚ�?             "@        ������������������������       �                     �?        u       x                    ?@      �?              @        v       w                 �̌!@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@        {       �                   �R@H�5�E6�?�            Pt@       |       �                    �? �qm���?�            �p@        }       �                     @�nN@��?I            �_@       ~       �                     �? 7���B�?,            @T@               �                   �H@H%u��?             9@       ������������������������       �                     4@        �       �                 �DD@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     L@        �       �                    �?X�<ݚ�?            �F@        ������������������������       �                     @        �       �                 ���7@�\��N��?             C@        �       �                    �?���N8�?             5@       �       �                   �/@�	j*D�?             *@        ������������������������       �                      @        �       �                    �?"pc�
�?             &@       ������������������������       �                     @        �       �                 @3�2@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �/@      �?              @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 X��@@�t����?             1@       ������������������������       �        	             *@        �       �                   @D@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?��|.V�?^             b@        �       �                    �?��
ц��?             :@        �       �                 �|�;@      �?	             ,@        ������������������������       �                     @        �       �                   �@@�z�G��?             $@        ������������������������       �                     @        �       �                   �J@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                 �|Y>@�q�q�?	             (@       �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                    *@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��&�F"�?L            �]@       �       �                    R@�'�`d�?C            �X@       �       �                    �?�����?B            �X@        �       �                 �|�2@      �?              @       ������������������������       �                     @        �       �                   `3@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �J@z�G�z�?=            �V@       �       �                   @I@�6i����?6            �S@       �       �                     �?6��f�?4            @S@        �       �                   �;@�t����?             A@        ������������������������       �                     �?        �       �                   �>@���!pc�?            �@@        �       �                 03:@և���X�?
             ,@        ������������������������       �                     @        �       �                 03k:@���!pc�?             &@        ������������������������       �                     �?        �       �                 �|Y=@�z�G��?             $@        ������������������������       �                     �?        �       �                   @G@�<ݚ�?             "@       �       �                 `fF<@����X�?             @       �       �                 �|�?@���Q��?             @        ������������������������       �                     �?        �       �                   �C@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @B@�}�+r��?             3@        ������������������������       �                      @        �       �                  x#J@�C��2(�?             &@        ������������������������       �                     @        �       �                    F@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 0�H@(L���?            �E@       �       �                    !@�X�<ݺ?             B@        �       �                   l@@����X�?             @       �       �                     @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     =@        �       �                 ��?P@և���X�?             @       �       �                    ;@z�G�z�?             @        ������������������������       �                     @        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        �       �                    $@�G�z��?	             4@       �       �                 pf�C@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                      @        �       �                   @E@�{��?��?&             K@       �       �                    �?���H��?             E@       �       �                    �?XB���?             =@       ������������������������       �                     ,@        �       �                    �?��S�ۿ?
             .@       ������������������������       �                     *@        �       �                 Ъ�c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�	j*D�?
             *@       �       �                    �?���|���?             &@       �       �                    �?����X�?             @       �       �                 X�,@@      �?             @       �       �                 �|Y;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �w|c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �̾w@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �                           �?      �?             (@       �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @                                 �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������KY� ��?iM���{�?���H	�?�T�/���?              �?q;x���?=�Y�?      �?        ��\V��?(፦ί�?0E>�S�?�u�)�Y�?d!Y�B�?ӛ���7�?              �?�?�������?F]t�E�?/�袋.�?�q�q�?9��8���?      �?              �?      �?              �?      �?                      �?              �?<<<<<<�?�?      �?        �l�w6��?AL� &W�?      �?        �������?�������?��{a�?a���{�?�������?�?۶m۶m�?�$I�$I�?      �?                      �?      �?        %I�$I��?�m۶m��?      �?      �?�$I�$I�?۶m۶m�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?        sƜ1g��?4�9c��?Ł�@q��?��u�:~�?;�;��?b'vb'v�?(�����?�k(���?              �?      �?      �?              �?      �?        e�M6�d�?6�d�M6�?      �?        I�$I�$�?n۶m۶�?333333�?�������?              �?�E]t��?]t�E]�?6��P^C�?(������?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?              �?      �?              �?      �?                      �?              �?|���?|���?�����?������?      �?      �?�m۶m��?�$I�$I�?              �?      �?        /�����?����X�?      �?        \��[���?�i�i�?ffffff�?�������?�q�q�?�q�q�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        6��P^C�?(������?              �?�������?UUUUUU�?�������?333333�?      �?                      �?�N��N��?ى�؉��?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?              �?        Y�Cc�?9/���?�m۶m��?�$I�$I�?      �?                      �?>��=���?��?      �?        �������?�?b�2�tk�?�����H�?      �?        �؉�؉�?;�;��?;�;��?;�;��?      �?      �?      �?        ��[��[�?�A�A�?      �?        �������?�������?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        9��8���?�q�q�?              �?      �?      �?�������?�������?      �?                      �?      �?              �?        �t|��?�������?	��3���?��f,�?�u]�u]�?��(��(�?h/�����?	�%����?���Q��?)\���(�?              �?333333�?�������?      �?                      �?              �?�q�q�?r�q��?              �?y�5���?�5��P�?��y��y�?�a�a�?;�;��?vb'vb'�?      �?        F]t�E�?/�袋.�?              �?�������?333333�?              �?      �?              �?      �?      �?      �?              �?      �?                      �?<<<<<<�?�?      �?              �?      �?              �?      �?        Q�k%��?^�(ٵ��?�;�;�?�؉�؉�?      �?      �?              �?ffffff�?333333�?      �?              �?      �?              �?      �?        �������?�������?UUUUUU�?�������?              �?      �?      �?              �?      �?              �?        8��7���?�k"�k"�?6�d�M6�?'�l��&�?^N��)x�?����X�?      �?      �?      �?              �?      �?      �?                      �?�������?�������?kq�w��?T:�g *�?g�'�Y�?�cj`��?�������?�������?              �?F]t�E�?t�E]t�?۶m۶m�?�$I�$I�?      �?        t�E]t�?F]t�E�?              �?333333�?ffffff�?      �?        �q�q�?9��8���?�$I�$I�?�m۶m��?�������?333333�?      �?              �?      �?              �?      �?      �?              �?              �?�5��P�?(�����?      �?        ]t�E�?F]t�E�?      �?        �������?UUUUUU�?              �?      �?        ⎸#��?w�qG��?��8��8�?�q�q�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ۶m۶m�?�$I�$I�?�������?�������?              �?      �?      �?      �?                      �?      �?                      �?      �?                      �?�������?�������?      �?      �?              �?      �?              �?        /�����?���^B{�?��y��y�?�0�0�?�{a���?GX�i���?              �?�?�������?              �?      �?      �?      �?                      �?;�;��?vb'vb'�?F]t�E�?]t�E]�?�$I�$I�?�m۶m��?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?              �?      �?      �?�m۶m��?�$I�$I�?              �?      �?        �������?�������?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�޵#hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                     @"��p�?�           8�@               c                  x#J@����>��?�            ps@              
                   �2@F�TȲ�?�            �i@               	                    �? �Cc}�?             <@                                  �1@���Q��?             @                                   3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@               ^                   �K@(����7�?q            @f@              W                   �G@,�Ѡ���?f            �d@              N                 �T�@@�L�w��?Y            �a@                                  �?�Cc}h,�?I             \@                                 s�,@�t����?             1@        ������������������������       �                     @                                    �?�q�q�?	             (@                                �>@      �?              @                                  B@�q�q�?             @                                Y>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @               1                    �?p�ݯ��?=            �W@               0                    :@�r����?             >@              /                    �?�J�4�?             9@                                  �'@r�q��?             8@        ������������������������       �                     @        !       (                    1@z�G�z�?             4@        "       #                    :@r�q��?             (@        ������������������������       �                     �?        $       %                   �A@�C��2(�?             &@       ������������������������       �                     @        &       '                    D@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        )       ,                   �7@      �?              @        *       +                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        -       .                   @B@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        2       3                    :@��ɉ�?)            @P@        ������������������������       �        
             0@        4       ?                     �?Jm_!'1�?            �H@        5       6                    <@���Q��?
             .@        ������������������������       �                      @        7       >                   @>@�	j*D�?	             *@       8       9                 ��:@ףp=
�?             $@        ������������������������       �                     @        :       =                 `f�;@z�G�z�?             @        ;       <                 �|�?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        @       A                   �@@l��\��?             A@        ������������������������       �        	             ,@        B       E                   @A@R���Q�?             4@        C       D                    1@      �?             @        ������������������������       �                      @        ������������������������       �                      @        F       M                    �?      �?	             0@       G       L                    ,@�8��8��?             (@        H       I                   �'@z�G�z�?             @        ������������������������       �                      @        J       K                   �C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        O       P                   �8@؇���X�?             <@        ������������������������       �                     @        Q       V                    �?`2U0*��?             9@       R       U                   �B@���N8�?             5@        S       T                 �|�<@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             .@        ������������������������       �                     @        X       Y                    �?�q�q�?             8@       ������������������������       �                     .@        Z       ]                   �I@�����H�?             "@        [       \                     �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        _       b                     �?@4և���?             ,@       `       a                   �R@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        d       �                    @���N8�?B            @Z@       e       f                    �?��[�8��?A            �Y@       ������������������������       �        (             P@        g       p                 ��4M@D�n�3�?             C@        h       i                    �?����X�?             @        ������������������������       �                      @        j       k                 `�iJ@���Q��?             @        ������������������������       �                     �?        l       m                    7@      �?             @        ������������������������       �                     �?        n       o                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        q       �                   @I@f���M�?             ?@       r       u                  �}S@
j*D>�?             :@        s       t                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        v       �                    �?�q�q�?             5@       w       �                    �?     ��?             0@       x                        @��v@�q�q�?             .@       y       ~                    �?�θ�?             *@       z       {                   @B@�q�q�?             "@        ������������������������       �                     @        |       }                   �H@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|�0@���Q��?             @        ������������������������       �                     �?        �       �                   �G@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�-���?�             y@        �       �                    �?�\��N��?C            �\@       �       �                    �?����S��?#             M@       �       �                   �-@     ��?             @@        �       �                   �,@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�9@@4և���?             <@        ������������������������       �                     @        �       �                    �?���}<S�?             7@        �       �                 ��%@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���@���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        �       �                   �@��
ц��?             :@        ������������������������       �                      @        �       �                 �|�=@�<ݚ�?
             2@       �       �                  �#@$�q-�?             *@       ������������������������       �                     &@        �       �                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   &@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �̼6@������?              L@        �       �                    �?���>4��?             <@        �       �                    &@�θ�?             *@        ������������������������       �                      @        �       �                 �|Y=@�C��2(�?             &@        �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �&@z�G�z�?             .@        �       �                 03c"@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�C��2(�?             &@       �       �                 pf�0@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��T?@؇���X�?             <@        ������������������������       �        	             .@        �       �                 ��p@@�	j*D�?	             *@        ������������������������       �                     @        ������������������������       �                     "@        �       �                    @8�Z$���?�            �q@        �       �                    �?�q�q�?             (@       �       �                 �Q��?      �?              @        ������������������������       �                      @        �       �                 ��|2@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?,�:\���?�             q@        �       �                 �|Y=@�q�q�?            �C@        �       �                   @@X�Cc�?
             ,@        �       �                   �5@�q�q�?             @        �       �                 �{@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    7@      �?              @        ������������������������       �                     @        �       �                   �;@z�G�z�?             @       �       �                 �0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�J�4�?             9@       �       �                 �|�=@���7�?             6@        �       �                 ���@�C��2(�?             &@        ������������������������       �                     @        �       �                 p&�@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        �                       �|�=@�;t~y�?�            `m@       �                       �T�I@t��ճC�?p             f@       �       �                    �?�}�+r��?m            `e@        ������������������������       �                     <@        �                          �?�'g�2�?^            �a@       �       �                 �?�@Du9iH��?U             `@       �       �                 �?$@��pBI�?/            @R@       �       �                    7@������?            �D@       ������������������������       �                     5@        �       �                 �&b@ףp=
�?             4@        ������������������������       �                     $@        �       �                 ���@z�G�z�?             $@        ������������������������       �                     �?        �       �                 �|�;@�����H�?             "@        ������������������������       �                     @        �       �                 pf�@r�q��?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @@        �       �                 @3�@      �?&             L@        �       �                   �4@      �?              @        ������������������������       �      �?             @        ������������������������       �                     @        �       �                   �3@�8��8��?!             H@        �       �                   �1@����X�?             @        ������������������������       �                     @        �       �                   �2@      �?             @        ������������������������       �                     �?        �       �                 `�8"@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        �       �                 ���"@������?            �D@       ������������������������       �                     6@        �                       `�X#@�KM�]�?             3@        �       �                   �<@���Q��?             @        ������������������������       �                      @        �                        �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �        	             ,@                              �|�;@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                                @@@$gv&��?$            �M@                                �>@b�2�tk�?
             2@        	      
                �̌!@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                �?@��
ц��?             *@        ������������������������       �                      @                                �@���|���?             &@        ������������������������       �                     @                              d�6@@և���X�?             @                             �?�@�q�q�?             @        ������������������������       �                     �?                              ��I @���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?                              @3�@��Y��]�?            �D@                              �?�@�X�<ݺ?             2@       ������������������������       �        
             1@        ������������������������       �                     �?        ������������������������       �                     7@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������J54v��?l�����?��f�?t�����?4��~���?�E|���?۶m۶m�?%I�$I��?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?<��x��?�9�as�?�JԮD��?%jW�v%�?|�W|�W�?uPuP�?%I�$I��?�m۶m��?�������?�������?              �?�������?�������?      �?      �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?                      �?      �?      �?              �?      �?        ^Cy�5�?Cy�5��?�?�������?{�G�z�?�z�G��?UUUUUU�?�������?              �?�������?�������?UUUUUU�?�������?      �?        F]t�E�?]t�E�?              �?�������?�������?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?                      �?              �?�����?�����?      �?        ����X�?������?333333�?�������?              �?vb'vb'�?;�;��?�������?�������?      �?        �������?�������?      �?      �?      �?                      �?      �?                      �?------�?�������?      �?        333333�?333333�?      �?      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ۶m۶m�?�$I�$I�?              �?���Q��?{�G�z�?��y��y�?�a�a�?�������?UUUUUU�?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?              �?�q�q�?�q�q�?      �?      �?              �?      �?              �?        n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?        ��y��y�?�a�a�?�������?�?              �?l(�����?(������?�$I�$I�?�m۶m��?              �?�������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��RJ)��?��Zk���?b'vb'v�?;�;��?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?ى�؉��?�؉�؉�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?      �?        333333�?�������?              �?      �?      �?      �?                      �?      �?              �?        �G�z��?�p=
ף�?�5��P�?y�5���?O#,�4��?X�i���?      �?      �?      �?      �?              �?      �?        �$I�$I�?n۶m۶�?              �?d!Y�B�?ӛ���7�?      �?      �?              �?      �?        �a�a�?��y��y�?      �?                      �?�;�;�?�؉�؉�?              �?9��8���?�q�q�?�؉�؉�?;�;��?      �?              �?      �?              �?      �?        �������?333333�?      �?                      �?I�$I�$�?n۶m۶�?n۶m۶�?I�$I�$�?ى�؉��?�؉�؉�?              �?]t�E�?F]t�E�?�������?�������?      �?                      �?      �?        �������?�������?      �?      �?              �?      �?        F]t�E�?]t�E�?UUUUUU�?�������?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?        vb'vb'�?;�;��?              �?      �?        ;�;��?;�;��?�������?�������?      �?      �?              �?�������?UUUUUU�?              �?      �?                      �?��ǭ�?ȭ�;�H�?UUUUUU�?UUUUUU�?�m۶m��?%I�$I��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?�z�G��?{�G�z�?�.�袋�?F]t�E�?]t�E�?F]t�E�?      �?        �������?UUUUUU�?�������?�������?      �?              �?                      �?Y�C�^��?5���	%�?�E]t��?t�E]t�?�5��P�?(�����?      �?        $T�ik��?�^���?qG�w��?w�qGܱ?���Ǐ�?����?p>�cp�?������?      �?        �������?�������?      �?        �������?�������?              �?�q�q�?�q�q�?      �?        �������?UUUUUU�?      �?              �?      �?      �?              �?      �?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?        p>�cp�?������?      �?        �k(���?(�����?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �������?333333�?              �?      �?        [4��}�?��/���?9��8���?�8��8��?�������?�������?      �?                      �?�؉�؉�?�;�;�?      �?        F]t�E�?]t�E]�?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?      �?      �?                      �?8��18�?������?��8��8�?�q�q�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�G�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM!hjh))��}�(h,h/h0M!��h2h3h4hph<�h=Kub������       6                   �1@�t����?�           8�@               #                 03�;@�X���?@             \@                                  /@�������?%             Q@                               ��-@��0{9�?            �G@        ������������������������       �        
             6@               	                    �? �o_��?             9@                                ��3@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        
                            @��s����?             5@       ������������������������       �                     &@                                   �?���Q��?             $@                                ��|2@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               "                    �?�G��l��?             5@                                 �0@�G�z��?             4@                                �̌!@      �?              @                                  �?r�q��?             @        ������������������������       �                     @                                pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                   �?�q�q�?             (@                                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                !                 ��)#@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        $       1                    )@�zv�X�?             F@       %       *                     @�E��ӭ�?             B@        &       )                    @���!pc�?             &@       '       (                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        +       0                    @HP�s��?             9@        ,       -                    �?�<ݚ�?             "@        ������������������������       �                     @        .       /                 ���A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             0@        2       5                 ���I@      �?              @        3       4                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        7       �                   �(@���\˾�?           ��@        8       W                    �?f?�ϼ��?�            `p@        9       J                    �?ٜSu��?,            @Q@        :       A                 �|Y=@      �?             B@        ;       @                   �<@���|���?             &@       <       ?                   �6@      �?              @        =       >                 ��y@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        B       C                    �?HP�s��?             9@        ������������������������       �                     �?        D       I                 �|�=@ �q�q�?             8@       E       F                 ���@�X�<ݺ?
             2@        ������������������������       �                     @        G       H                   @@�8��8��?             (@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     @        K       R                    �?:ɨ��?            �@@        L       Q                    �?X�Cc�?
             ,@       M       N                 �|�9@ףp=
�?	             $@        ������������������������       �                      @        O       P                  ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        S       V                 X��A@�}�+r��?             3@       T       U                 �Y�@��S�ۿ?
             .@        ������������������������       �                     @        ������������������������       ��8��8��?             (@        ������������������������       �                     @        X       Y                 ���@�ը
q��?             h@        ������������������������       �                     6@        Z       s                    �?^<����?p            `e@        [       p                 �|�?@|��?���?             ;@       \       ]                     @և���X�?             5@        ������������������������       �                     �?        ^       c                   �@���Q��?             4@        _       `                 ���@r�q��?             @        ������������������������       �                     @        a       b                    4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        d       m                    �?d}h���?
             ,@       e       f                   �3@z�G�z�?             $@        ������������������������       �                     �?        g       l                 @3�@�����H�?             "@        h       i                 �?�@      �?             @        ������������������������       �                      @        j       k                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        n       o                   �#@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        q       r                   �J@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        t       u                 ���@���Hx�?[             b@        ������������������������       �                      @        v       �                   �<@@�j;��?Z            �a@        w       |                     @0�,���?+            �P@        x       y                   �2@      �?              @        ������������������������       �                     @        z       {                   �5@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        }       ~                 �?�@P����?&            �M@       ������������������������       �                     B@               �                 0S5 @�nkK�?             7@        �       �                   �3@      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �        
             .@        �       �                     @�r����?/            �R@        ������������������������       �                     (@        �       �                   @@@��d��?)            �O@       �       �                 �|Y>@      �?             B@       �       �                 ���"@      �?             8@       �       �                 �|Y=@���}<S�?             7@        ������������������������       �                     @        �       �                  sW@�KM�]�?             3@        �       �                 ��,@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             (@        ������������������������       �                     �?        �       �                   �?@      �?             (@        ������������������������       �                     �?        �       �                   �@�eP*L��?             &@        ������������������������       �                     @        �       �                 �?�@      �?              @        ������������������������       �                     �?        �       �                 ��I @����X�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                 @3�@ 7���B�?             ;@       �       �                 �?�@�8��8��?
             (@       ������������������������       �                     $@        ������������������������       �      �?              @        ������������������������       �                     .@        �       �                 `fK@8�lC(��?�            u@       �       �                    �?n�.P���?�             o@        �       �                    @6�"W�u�?A            �Y@       �       �                    �?��8����?<             X@       �       �                 ��0@�qM�R��?(            �P@        ������������������������       �                     9@        �       �                   �3@؇���X�?             E@        �       �                 03�0@և���X�?             @       �       �                 �|�;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                     �? >�֕�?            �A@        �       �                    �?      �?             0@        �       �                   �H@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             3@        �       �                    �?>���Rp�?             =@       �       �                     @�E��ӭ�?             2@        ������������������������       �                     $@        �       �                   �>@      �?              @       �       �                   �6@����X�?             @        ������������������������       �                      @        �       �                 �A7@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|Y=@"pc�
�?             &@       ������������������������       �                      @        �       �                 �|Y?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �C@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?д>��C�?Z             b@       �       �                     �?�0*��?N            �_@        �       �                    �?���dQ'�?#            �L@        �       �                  Y>@�8��8��?             (@        �       �                 ���=@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�<@k��9�?            �F@        �       �                    7@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        �       �                  i?@      �?             @@       �       �                   @=@b�2�tk�?             2@       �       �                 `f�;@������?	             .@       �       �                 `fF:@�q�q�?             (@        ������������������������       �                      @        �       �                   �K@���Q��?             $@       �       �                 �|�?@և���X�?             @        ������������������������       �                      @        �       �                   �C@z�G�z�?             @        ������������������������       �                      @        �       �                   @G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                  x#J@@4և���?
             ,@       ������������������������       �                     $@        �       �                   �C@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �*@ >�֕�?+            �Q@        �       �                    �?"pc�
�?             6@        ������������������������       �                     �?        �       �                 �|Y<@��s����?             5@        ������������������������       �                     @        �       �                 `f�)@������?	             .@        ������������������������       �                     �?        �       �                 �|�=@����X�?             ,@        ������������������������       �                      @        �       �                    @@r�q��?             (@        ������������������������       �                     @        �       �                   �F@      �?              @       �       �                   @D@���Q��?             @       �       �                   @B@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     H@        �       �                   �6@�X�<ݺ?             2@        ������������������������       �                     �?        ������������������������       �                     1@        �       
                �|�=@\{��)x�?9            @V@        �       �                 @3[Q@և���X�?            �A@        �       �                    �?؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @               	                    �?�ՙ/�?             5@                              �k@      �?             0@                                �?�z�G��?             $@       ������������������������       �                     @                               �}S@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                 5@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                               `D�c@�{��?��?#             K@                             �UcV@      �?             F@                                �?8�Z$���?             :@        ������������������������       �                     ,@                                 �?�q�q�?             (@                                  @�����H�?             "@                                �?؇���X�?             @       ������������������������       �                     @                              03�M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?b�2�tk�?             2@       ������������������������       �                      @                                 �?�z�G��?             $@                                �G@���Q��?             @        ������������������������       �                     �?                                 �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �*       h�h))��}�(h,h/h0M!KK��h2h3h4hVh<�h=Kub������������G�+J>�?r%�k���?n۶m۶�?I�$I�$�?�������?�������?L� &W�?m�w6�;�?              �?�Q����?
ףp=
�?      �?      �?      �?                      �?�a�a�?z��y���?              �?�������?333333�?۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?1�0��?��y��y�?�������?�������?      �?      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?��.���?�袋.��?�q�q�?r�q��?t�E]t�?F]t�E�?      �?      �?              �?      �?                      �?q=
ףp�?{�G�z�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?��@?�?�:z�~��?�]�WqB�?ˈ>�:��?s��\;0�?%~F���?      �?      �?F]t�E�?]t�E]�?      �?      �?�������?�������?      �?                      �?      �?                      �?q=
ףp�?{�G�z�?              �?�������?UUUUUU�?��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?              �?        N6�d�M�?e�M6�d�?�m۶m��?%I�$I��?�������?�������?              �?      �?      �?      �?                      �?      �?        �5��P�?(�����?�������?�?      �?        UUUUUU�?UUUUUU�?      �?        ��
��[�?����?      �?        *������?XOa=���?	�%����?{	�%���?�$I�$I�?۶m۶m�?              �?333333�?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?I�$I�$�?۶m۶m�?�������?�������?              �?�q�q�?�q�q�?      �?      �?      �?              �?      �?      �?                      �?      �?              �?      �?              �?      �?        UUUUUU�?�������?              �?      �?        9��8���?9��8��?              �?w�'�K�?H���@��?Ez�rv�?g��1��?      �?      �?      �?        �������?�������?      �?      �?      �?        �V'u�?'u_[�?      �?        �Mozӛ�?d!Y�B�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?        �������?�?      �?        ��뺮��?EQEQ�?      �?      �?      �?      �?ӛ���7�?d!Y�B�?      �?        �k(���?(�����?�m۶m��?�$I�$I�?      �?                      �?      �?                      �?      �?      �?              �?t�E]t�?]t�E�?              �?      �?      �?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?        	�%����?h/�����?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        ��)�8%�?k�cm�?�9�s��?c�1�c�?#>�Tr^�?w��jch�?UUUUUU�?�������?���@��?�n�Wc"�?              �?�$I�$I�?۶m۶m�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?        �A�A�?��+��+�?      �?      �?F]t�E�?/�袋.�?              �?      �?                      �?              �?GX�i���?�i��F�?r�q��?�q�q�?              �?      �?      �?�m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?                      �?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?�m۶m��?�$I�$I�?              �?      �?        a���{�?|a���?}>�����?��`0�?ZLg1���?Lg1��t�?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?        �'}�'}�?[�[��?;�;��?;�;��?      �?                      �?      �?      �?�8��8��?9��8���?wwwwww�?�?UUUUUU�?UUUUUU�?      �?        333333�?�������?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?n۶m۶�?�$I�$I�?      �?              �?      �?      �?                      �?��+��+�?�A�A�?/�袋.�?F]t�E�?      �?        z��y���?�a�a�?      �?        wwwwww�?�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ��8��8�?�q�q�?              �?      �?        +Y�JV��?jS��Ԧ�?۶m۶m�?�$I�$I�?�$I�$I�?۶m۶m�?              �?      �?        �<��<��?�a�a�?      �?      �?333333�?ffffff�?              �?      �?      �?              �?      �?        �������?UUUUUU�?              �?      �?              �?        /�����?���^B{�?      �?      �?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?      �?        9��8���?�8��8��?              �?ffffff�?333333�?�������?333333�?      �?              �?      �?      �?                      �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���JhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       J                    �?���;+"�?�           8�@               3                    �?և���X�?U            @c@                                  �?@lܯ ��?@            �]@                                0Cd=@�NW���?            �J@                                    �?����X�?	             ,@        ������������������������       �                      @                                �|�<@r�q��?             (@                                 �-@ףp=
�?             $@        	       
                   �+@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                ��%@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �C@                                �|Y=@r٣����?&            �P@                                0C�<@�\��N��?             3@                               �&�)@X�Cc�?	             ,@                               ��=@����X�?             @                                  5@�q�q�?             @        ������������������������       �                     �?                                  �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                �U�X@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?               2                 p�w@��0{9�?            �G@               1                   `E@�C��2(�?             F@       !       0                   �B@(N:!���?            �A@       "       '                     �?l��\��?             A@        #       &                 ��2>@r�q��?             (@        $       %                 ���<@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        (       )                 ���@���7�?             6@        ������������������������       �                     "@        *       +                     @$�q-�?	             *@        ������������������������       �                      @        ,       /                 �|Y?@�C��2(�?             &@       -       .                   @@؇���X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        4       ?                     �?^������?            �A@        5       <                    �?     ��?	             0@       6       7                    �?��
ц��?             *@        ������������������������       �                     @        8       9                 ��UO@      �?              @        ������������������������       �                     @        :       ;                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        =       >                    C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        @       A                 ���,@�S����?             3@        ������������������������       �                     @        B       E                    �?     ��?
             0@        C       D                 `f�=@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        F       I                 `�@1@      �?              @        G       H                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        K       �                     @��6��?V           h�@        L       e                    �?\�>�6��?�            `o@        M       `                 ���a@ЮN
��?A            @\@       N       _                    �?@9G��?:            �X@       O       X                   �;@`Jj��?$             O@        P       Q                     �?      �?             (@        ������������������������       �                     @        R       S                   �5@      �?              @        ������������������������       �                     @        T       W                   �9@���Q��?             @       U       V                   �3@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        Y       Z                  ��9@p���?             I@        ������������������������       �                     9@        [       \                   �E@`2U0*��?             9@       ������������������������       �                     4@        ]       ^                 `fF:@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     B@        a       d                 Ъ�c@�r����?             .@        b       c                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        f       g                    $@��<b���?V            @a@        ������������������������       �                     @        h       �                     �?|�-蝉�?S            �`@        i       j                    �?N{�T6�?!            �K@        ������������������������       �                     �?        k       �                    �?b�2�tk�?              K@       l       �                 ��9L@���H.�?             I@       m       ~                  i?@F�����?            �F@       n       }                   �L@��
ц��?             :@       o       |                   `G@���|���?             6@       p       {                   �B@��.k���?
             1@       q       r                 ��I*@      �?             (@        ������������������������       �                     �?        s       z                 `f�<@"pc�
�?             &@       t       u                 �|�<@      �?              @        ������������������������       �                     @        v       w                 03k:@���Q��?             @        ������������������������       �                      @        x       y                 �|�?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               �                   �C@�S����?             3@       �       �                 �|�<@�8��8��?             (@        �       �                   �7@z�G�z�?             @        ������������������������       �                     �?        �       �                 `f�D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @F@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @C@z�G�z�?             @        ������������������������       �                     @        �       �                 XfZX@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�7��?2            �S@       �       �                   �E@�}�+r��?0             S@       �       �                   @D@ ,��-�?&            �M@       �       �                    @�1�`jg�?#            �K@        ������������������������       �                     $@        �       �                    1@��S�ۿ?            �F@       �       �                   �(@�#-���?            �A@       �       �                    5@�X�<ݺ?             2@        �       �                    &@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     (@        �       �                 �|�<@�t����?             1@        ������������������������       �                     @        �       �                 �|�=@z�G�z�?             $@        ������������������������       �                     �?        �       �                   �A@�����H�?             "@       �       �                    @@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    4@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �        
             1@        ������������������������       �                      @        �       �                 ���@������?�             s@        ������������������������       �                     5@        �                         @1@�ț��*�?�            �q@       �       �                   �1@���{��?�            `k@        �       �                    �?�}�+r��?             3@       ������������������������       �                     &@        �       �                    �?      �?              @        �       �                 pf�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?H.�!���?             i@        �       �                   �7@      �?             D@        ������������������������       �                     @        �       �                    �?4�B��?            �B@       �       �                    �?ҳ�wY;�?             A@        ������������������������       �                     &@        �       �                 �|Y;@�nkK�?             7@        ������������������������       �                     �?        �       �                 ��(@���7�?             6@       �       �                 ���@�X�<ݺ?
             2@        ������������������������       �                      @        ������������������������       �      �?             0@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��Q���?g             d@        �       �                   �C@l��[B��?             =@       �       �                    �?
j*D>�?             :@       �       �                 pf�@� �	��?             9@        ������������������������       �                     @        �       �                    �?�G��l��?             5@       �       �                 ��&@��.k���?             1@       �       �                   �3@�	j*D�?             *@        ������������������������       �                     @        �       �                   �@ףp=
�?             $@        �       �                 �&B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @C@A5Xo�?T            ``@       �       �                    �?�t`�4 �?M            �^@       �       �                   �:@�C��2(�?L            @^@        �       �                 ���@ 7���B�?"             K@        ������������������������       �                     �?        �       �                 �?�@�O4R���?!            �J@       ������������������������       �                    �@@        �       �                 @3�@P���Q�?             4@        �       �                   �4@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     0@        �       �                   �;@��v����?*            �P@        �       �                 �� @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �Yu@�����?(            �O@        �       �                 P��@�q�q�?             (@        ������������������������       �                     @        �       �                 �&B@X�<ݚ�?             "@       �       �                 �|Y>@և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y=@`'�J�?!            �I@        �       �                 ���"@      �?              @       ������������������������       �                     @        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�@ qP��B�?            �E@        �       �                    ?@��S�ۿ?             .@       ������������������������       �        	             (@        ������������������������       ��q�q�?             @        ������������������������       �                     <@        ������������������������       �                     �?        �                          �?�q�q�?             "@       �                        �?�@      �?              @        ������������������������       �                      @                              @3�@      �?             @        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?                              �T�I@6YE�t�?'            �P@                             ��p@@�?�P�a�?$             N@                             ��T?@fP*L��?             F@                                �?��(\���?             D@       	                         �?�S����?             3@        
                      X�,A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                              �|Y>@      �?
             0@       ������������������������       �                     *@                                 C@�q�q�?             @                             03C3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     @        ������������������������       �        
             0@                                 �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������D�#{��?x��	��?۶m۶m�?�$I�$I�?��
��
�?1�z1�z�?�x+�R�?萚`���?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?                      �?>���>�?|���?y�5���?�5��P�?%I�$I��?�m۶m��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        �������?�������?              �?      �?        m�w6�;�?L� &W�?]t�E�?F]t�E�?|�W|�W�?�A�A�?------�?�������?�������?UUUUUU�?333333�?�������?      �?                      �?      �?        �.�袋�?F]t�E�?      �?        �؉�؉�?;�;��?      �?        ]t�E�?F]t�E�?۶m۶m�?�$I�$I�?      �?      �?      �?              �?                      �?      �?                      �?_�_��?uPuP�?      �?      �?�;�;�?�؉�؉�?              �?      �?      �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ^Cy�5�?(������?              �?      �?      �?      �?      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?	�L])��?�}fE��?�Tw�V�?�UD�Tw�?4��A�/�?m���M�?9/���?������?�B!��?���{��?      �?      �?              �?      �?      �?              �?333333�?�������?      �?      �?      �?                      �?      �?        {�G�z�?\���(\�?              �?{�G�z�?���Q��?              �?�������?�������?      �?                      �?              �?�?�������?      �?      �?              �?      �?                      �?��,d!�?��Moz��?              �?	&��?���f�?�S�<%��?pX���o�?      �?        �8��8��?9��8���?���(\��?�z�G��?�>�>��?؂-؂-�?�؉�؉�?�;�;�?F]t�E�?]t�E]�?�?�������?      �?      �?      �?        F]t�E�?/�袋.�?      �?      �?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?      �?        (������?^Cy�5�?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?              �?        �m۶m��?�$I�$I�?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?      �?        ��[��[�?�A�A�?�5��P�?(�����?[4���?'u_[�?A��)A�?�־a�?      �?        �������?�?�A�A�?_�_�?��8��8�?�q�q�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        <<<<<<�?�?      �?        �������?�������?              �?�q�q�?�q�q�?�������?�������?      �?              �?      �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?              �?        xxxxxx�?�?      �?        �~�-q��?�a�+�?o3����?�!��d�?(�����?�5��P�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�(\����?)\���(�?      �?      �?              �?�Y7�"��?L�Ϻ��?�������?�������?              �?�Mozӛ�?d!Y�B�?      �?        �.�袋�?F]t�E�?��8��8�?�q�q�?      �?              �?      �?      �?              �?        333333�?333333�?GX�i���?���=��?;�;��?b'vb'v�?)\���(�?�Q����?              �?1�0��?��y��y�?�������?�?vb'vb'�?;�;��?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?      �?              �?      �?                      �?      �?        ��℔�?#����[�?~�K�`�?�����?]t�E�?F]t�E�?	�%����?h/�����?              �?:�&oe�?�x+�R�?      �?        ffffff�?�������?      �?      �?      �?      �?      �?              �?        5&����?*g��1�?      �?      �?      �?                      �?=��<���?�a�a�?UUUUUU�?UUUUUU�?      �?        r�q��?�q�q�?�$I�$I�?۶m۶m�?�������?333333�?      �?              �?      �?      �?                      �?�������?�?      �?      �?      �?              �?      �?      �?                      �?��}A�?�}A_З?�������?�?      �?        UUUUUU�?UUUUUU�?      �?              �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?      �?      �?              �?        '�l��&�?e�M6�d�?DDDDDD�?�����ݽ?颋.���?]t�E]�?�������?333333�?(������?^Cy�5�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?      �?              �?      �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�
HyhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0Kᅔh2h3h4hph<�h=Kub��������       X                    �?��ϙLq�?�           8�@               U                    @f��>���?�            �o@              >                 �|�=@D4�K�p�?�            �n@              =                 �̌R@���f+�?k            `e@              <                 @3[Q@2p�ZAJ�?a            �c@                                   @¦	^_�?_            `c@        ������������������������       �                     H@                                   �?�"��61�?@            �Z@        	                           �?>A�F<�?             C@        
                           @�n_Y�K�?             *@                               H�%@      �?             $@        ������������������������       �                     @                                  �@����X�?             @        ������������������������       �                     �?                                03�-@r�q��?             @                                 �-@      �?             @        ������������������������       �                      @                                  �0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                ���@HP�s��?             9@        ������������������������       �                      @        ������������������������       �                     7@                                   @��z4���?(            @Q@                                   �?�����H�?             "@                               @3�2@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                !                   �0@�0u��A�?"             N@        ������������������������       �                     (@        "       ;                 ��Y1@�q���?             H@       #       $                   �1@d�
��?             F@        ������������������������       �                     @        %       8                 �|�<@�Q����?             D@       &       7                   �;@���Q��?             >@       '       (                 pf�@�q�����?             9@        ������������������������       �                     @        )       6                    �?�ՙ/�?             5@       *       5                 pf� @     ��?             0@        +       0                 �&B@      �?              @        ,       -                    4@z�G�z�?             @        ������������������������       �                     @        .       /                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       2                 P�@�q�q�?             @        ������������������������       �                     �?        3       4                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        9       :                 pf&(@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             (@        ?       P                     @@݈g>h�?.             S@       @       M                   @L@ =[y��?(             Q@       A       B                     �?�]0��<�?#            �N@       ������������������������       �                     A@        C       L                   @F@�>����?             ;@       D       K                   �E@؇���X�?	             ,@       E       J                   @0@$�q-�?             *@       F       G                   �A@      �?              @       ������������������������       �                     @        H       I                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        N       O                   �L@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        Q       T                   @D@      �?              @        R       S                 03�1@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        V       W                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        Y       �                    �?��)�c{�?)           �|@        Z       q                 ��K.@H�U?B�?5            �T@        [       p                 �&�)@x�����?            �C@       \       o                 pF�#@r٣����?            �@@       ]       n                 �-!@     ��?             @@       ^       e                   @9@>���Rp�?             =@        _       `                 ���@      �?              @        ������������������������       �                      @        a       b                    �?      �?             @        ������������������������       �                      @        c       d                 ��}@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        f       g                 ���@�����?             5@        ������������������������       �                     "@        h       m                 �|�=@r�q��?	             (@       i       l                   @@�<ݚ�?             "@       j       k                 �|=@����X�?             @        ������������������������       �                      @        ������������������������       ����Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        r       �                    �?X��ʑ��?            �E@       s       x                 �|Y<@���Q��?             9@        t       w                 8��B@      �?              @        u       v                   �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        y       �                 xSQ@������?             1@       z       {                   @@@     ��?             0@        ������������������������       �                     @        |       �                 p�i@@�z�G��?             $@       }       �                  �>@      �?             @       ~                          �F@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                     @b�2�tk�?
             2@       �       �                     �?���|���?             &@       �       �                    �?���Q��?             $@       �       �                 ��UO@      �?             @        ������������������������       �                      @        �       �                 0��U@      �?             @        ������������������������       �                      @        �       �                   @E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �Q��?�C��2(�?�            `w@        ������������������������       �                     @        �       �                    #@�L���?�             w@        �       �                     @�q�q�?             5@        ������������������������       �                     @        �       �                    �?�<ݚ�?             2@        ������������������������       �                     @        �       �                 ���4@������?             .@        ������������������������       �                     @        ������������������������       �                     &@        �       �                 `fF:@��ϫ���?�            �u@       �       �                    �?����=O�?�             r@        �       �                   `3@XB���?             =@       ������������������������       �                     9@        �       �                 03�7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 @3�@�.^J��?�            Pp@        �       �                     @��X��?E             \@        ������������������������       �                     *@        �       �                    �?�C��2(�??            �X@       �       �                 �?�@�)���Y�?>            �X@       �       �                 ��L@��+��<�?8            �U@       ������������������������       �        !             I@        �       �                    ?@�8��8��?             B@       ������������������������       �                     >@        �       �                   �@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �A@      �?             (@       �       �                   �4@���Q��?             $@        ������������������������       ��q�q�?             @        �       �                   �:@����X�?             @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �3@@m����?a            �b@        �       �                   �2@P���Q�?             4@       ������������������������       �        
             *@        �       �                 0S5 @؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                     @�7�	|��?R             `@        �       �                 �|�=@ �Jj�G�?#            �K@        �       �                   �(@�}�+r��?             3@        ������������������������       �                     @        �       �                 �|Y=@�8��8��?	             (@       ������������������������       �                     $@        �       �                 `fv3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     B@        ������������������������       �        /            �R@        �       �                    R@F�4�Dj�?*            �M@       �       �                    �?д>��C�?)             M@       �       �                  i?@�<ݚ�?!            �F@        �       �                     �?X�<ݚ�?             2@       �       �                   @>@��.k���?             1@       �       �                 `fF<@X�Cc�?	             ,@       �       �                   �J@�q�q�?             (@       �       �                   @G@z�G�z�?             @        �       �                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �B@�>����?             ;@       ������������������������       �                     .@        �       �                   �E@r�q��?	             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     *@        ������������������������       �                     �?        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������Ӭ����?�X�>��?�������?�?S���.�?�W���?m%���V�?Im%����?Eg@(��?]z��k#�?�RJ)���?��Zk���?              �?��L�w��?9��/Ċ�?Cy�5��?������?ى�؉��?;�;��?      �?      �?              �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?      �?      �?              �?      �?              �?      �?              �?                      �?{�G�z�?q=
ףp�?      �?                      �?%~F���?̵s���?�q�q�?�q�q�?�$I�$I�?۶m۶m�?              �?      �?                      �?�������?�������?      �?        �������?�������?�.�袋�?�袋.��?              �?�������?ffffff�?333333�?�������?�p=
ף�?���Q��?              �?�<��<��?�a�a�?      �?      �?      �?      �?�������?�������?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?      �?        333333�?ffffff�?      �?                      �?      �?              �?                      �?Cy�5��?�P^Cy�?�������?�������?;ڼOqɠ?\2�h��?              �?h/�����?�Kh/��?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?�������?�������?              �?      �?              �?              �?      �?              �?      �?        Cy�5��?��k(��?�D�JԮ�?�v%jW��?��o��o�?�A�A�?>���>�?|���?      �?      �?�i��F�?GX�i���?      �?      �?              �?      �?      �?              �?      �?      �?      �?                      �?=��<���?�a�a�?      �?        �������?UUUUUU�?9��8���?�q�q�?�m۶m��?�$I�$I�?      �?        333333�?�������?      �?              �?              �?                      �?      �?        �}A_�?��}A�?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?xxxxxx�?�?      �?      �?      �?        ffffff�?333333�?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?9��8���?�8��8��?]t�E]�?F]t�E�?333333�?�������?      �?      �?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?              �?      �?              �?                      �?]t�E�?F]t�E�?              �?}���g�?L�Ϻ��?UUUUUU�?UUUUUU�?              �?9��8���?�q�q�?      �?        wwwwww�?�?              �?      �?        5kF ��?Y>���ް?U��K��?��RA�/�?GX�i���?�{a���?      �?              �?      �?              �?      �?        ��H���?��v��?۶m۶m�?%I�$I��?      �?        ]t�E�?F]t�E�?Dc}h��?������?�#�;��?w�qGܡ?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?333333�?�������?UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?        2�O
��?�3�=l}�?ffffff�?�������?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        ����?���?k߰�k�?��)A��?�5��P�?(�����?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?        ��/���?�A�I��?a���{�?|a���?9��8���?�q�q�?r�q��?�q�q�?�������?�?%I�$I��?�m۶m��?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?      �?              �?      �?      �?                      �?              �?      �?        �Kh/��?h/�����?      �?        �������?UUUUUU�?              �?      �?              �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���]hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       f                    �?�����?�           8�@               Q                    �?      �?�            �o@                                   @     ��?{             h@                               0Cd=@Xl���?E            �\@                                  �?�^����?%            �M@                                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        	                          �;@4��?�?!             J@        
                          �6@���!pc�?             &@       ������������������������       �                     @                                   8@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                ���&@������?            �D@                                  �J@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?                                   �?      �?             @@        ������������������������       �                     @                                  �E@XB���?             =@       ������������������������       �                     7@                                    �?r�q��?             @        ������������������������       �                     @                                  @F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �K@               .                 �̌@�e����?6            �S@               -                 X��B@�>4և��?             <@              &                    �?ȵHPS!�?             :@               %                 ���@��S�ۿ?             .@        !       "                 �|Y5@z�G�z�?             @        ������������������������       �                     �?        #       $                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        '       (                   �2@"pc�
�?             &@        ������������������������       �                     �?        )       ,                 pf�@ףp=
�?             $@        *       +                 �|Y:@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        /       6                    @z�):���?#             I@        0       1                    �?      �?              @        ������������������������       �                     @        2       3                    @z�G�z�?             @        ������������������������       �                      @        4       5                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        7       P                 �A7@�ՙ/�?             E@       8       K                 ��.@D�n�3�?             C@       9       <                    3@�q�q�?             >@        :       ;                   �-@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        =       >                    �?���y4F�?             3@        ������������������������       �                      @        ?       H                 ��&@������?             1@       @       G                 �|Y>@؇���X�?             ,@       A       B                   �9@$�q-�?
             *@       ������������������������       �                     $@        C       D                 �?�@�q�q�?             @        ������������������������       �                     �?        E       F                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        I       J                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        L       M                 03�1@      �?              @        ������������������������       �                     @        N       O                 `v�5@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        R       [                 03�;@���Q��?!             N@        S       T                     @H%u��?             9@       ������������������������       �                     .@        U       Z                 �|Y=@�z�G��?             $@       V       W                    �?      �?              @        ������������������������       �                     @        X       Y                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        \       ]                 ��T?@���Q��?            �A@        ������������������������       �                     (@        ^       a                     @�û��|�?             7@       _       `                    @�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        b       c                    @���!pc�?             &@        ������������������������       �                      @        d       e                    @�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        g       t                    $@"~��F��?(           �|@        h       m                   �;@�ՙ/�?             5@       i       l                    @$�q-�?	             *@        j       k                     @؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        n       o                    �?      �?              @        ������������������������       �                     @        p       s                    @      �?             @       q       r                 pf�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        u       �                     �?^	����?           `{@        v       �                  �>@�t����?=            �Y@        w       x                 `fF:@~�4_�g�?             F@        ������������������������       �                     $@        y       �                    �?�ʻ����?             A@       z       �                    @@���@M^�?             ?@        {       |                    <@�q�q�?             (@        ������������������������       �                     @        }       ~                   �<@�<ݚ�?             "@        ������������������������       �                     @               �                   @>@�q�q�?             @       �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �J@�d�����?
             3@       �       �                 `f�;@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        �       �                 `fF<@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @I@&y�X���?$             M@       �       �                    �?      �?             F@       �       �                    �?����>�?            �B@        �       �                 @�6M@�����?
             3@        ������������������������       �                     @        �       �                 @�pX@      �?             (@        �       �                   �9@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 X�,@@z�G�z�?             @        ������������������������       �                      @        �       �                 �Vs@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|Y<@�<ݚ�?             2@        ������������������������       �                      @        �       �                   @H@      �?             0@       �       �                 `f�K@��S�ۿ?
             .@       ������������������������       �                     $@        �       �                 03�M@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �B@؇���X�?             @       �       �                   �?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             ,@        �       �                 �?�@�Cc}h��?�             u@        �       �                    �?@ݚ)�?b             b@        �       �                   �6@ףp=
�?             >@        �       �                    �?      �?             @       �       �                 ��y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���@ ��WV�?             :@       ������������������������       �        	             ,@        �       �                 �|=@�8��8��?             (@        ������������������������       �                     @        �       �                 �|�=@      �?              @       �       �                   @@r�q��?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �?$@0�)AU��?M            �\@       �       �                    7@��
���?2            �R@        ������������������������       �                     5@        �       �                   �8@ 7���B�?&             K@        �       �                 `fF@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �? pƵHP�?$             J@        ������������������������       �                     4@        �       �                 pf�@      �?             @@       ������������������������       �                     <@        �       �                 �|�;@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                    �C@        �       �                 @3�@8��8���?z             h@        �       �                   �=@      �?             0@        ������������������������       �                     @        �       �                   �?@���!pc�?             &@        ������������������������       �                     @        �       �                   �A@և���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �      �?             @        �       �                   �4@�Ra����?r             f@        �       �                   �2@������?             ;@       �       �                     @�t����?             1@        ������������������������       �                     @        �       �                 pf� @8�Z$���?	             *@        �       �                    1@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?      �?             $@        ������������������������       �                     �?        �       �                     @X�<ݚ�?             "@        ������������������������       �      �?              @        �       �                 0S5 @և���X�?             @       �       �                   �3@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                      @        �                         @A@�
�@c�?_            �b@       �       �                 ��) @ܔQ|ӭ�?G            �[@        ������������������������       �                     9@        �       	                   �?,�"���?;            @U@       �       �                    �?�?�'�@�?5             S@        �       �                 ��$1@$�q-�?
             *@       ������������������������       �                      @        �       �                 м;4@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��y @؇���X�?+            �O@        ������������������������       �                      @        �       �                     @Xny��?*            �N@        �       �                 �|Y=@�����H�?             ;@        ������������������������       �        	             *@        �       �                 `fF)@d}h���?
             ,@        ������������������������       �                     @        �       �                 �|�=@���!pc�?             &@        ������������������������       �                      @        �       �                    @@�����H�?             "@        ������������������������       �                     @        �       �                    1@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        �                       ��C@�t����?             A@       �                          (@     ��?             @@       �                       ���"@؇���X�?             5@       �                          <@�IєX�?	             1@       �                          �:@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@                                �<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@                              �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        
                         �?�q�q�?             "@                                 @���Q��?             @        ������������������������       �                     �?                                 �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�����������������?��܍��?      �?      �?      �?     ��?��Gp�?��>���?W'u_�?u_[4�?�$I�$I�?�m۶m��?      �?                      �?ى�؉��?�N��N��?t�E]t�?F]t�E�?              �?      �?      �?      �?                      �?������?p>�cp�?�q�q�?�q�q�?              �?      �?              �?      �?              �?�{a���?GX�i���?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?�A�A�?�-��-��?�m۶m��?�$I�$I�?�؉�؉�?��N��N�?�?�������?�������?�������?              �?      �?      �?              �?      �?                      �?F]t�E�?/�袋.�?      �?        �������?�������?      �?      �?              �?      �?                      �?      �?        H�z�G�?q=
ףp�?      �?      �?              �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �<��<��?�a�a�?l(�����?(������?UUUUUU�?UUUUUU�?]t�E�?t�E]t�?      �?                      �?6��P^C�?(������?      �?        xxxxxx�?�?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?333333�?���Q��?)\���(�?              �?333333�?ffffff�?      �?      �?              �?      �?      �?              �?      �?              �?        333333�?�������?      �?        ��,d!�?8��Moz�?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?                      �?�A^%���?���j�1�?�a�a�?�<��<��?;�;��?�؉�؉�?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?      �?      �?              �?      �?      �?      �?              �?      �?              �?        [�lٲe�?�&M�4i�?�������?�������?/�袋.�?��.���?      �?        <<<<<<�?�������?�c�1��?�s�9��?�������?�������?              �?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?y�5���?Cy�5��?;�;��?�؉�؉�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ��FX��?�i��F�?      �?      �?�u�)�Y�?���L�?Q^Cy��?^Cy�5�?      �?              �?      �?�$I�$I�?�m۶m��?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?9��8���?�q�q�?              �?      �?      �?�������?�?      �?        �������?�������?              �?      �?                      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �m۶m��?I�$I�$�?9��8���?r�qǡ?�������?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        O��N���?;�;��?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?�������?UUUUUU�?�������?�������?      �?              �?        ��Gp�?p�}��?&�X�%�?O贁N�?      �?        	�%����?h/�����?      �?      �?              �?      �?        'vb'vb�?;�;��?      �?              �?      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?�������?      �?      �?      �?        t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?]t�E]�?]t�E�?B{	�%��?{	�%���?<<<<<<�?�?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?      �?              �?r�q��?�q�q�?      �?      �?�$I�$I�?۶m۶m�?�������?333333�?      �?      �?      �?              �?        �ַC5�?�IA��U�?8�}��7�?A��)A�?      �?        �?�������?������?y�5���?�؉�؉�?;�;��?      �?        �������?�������?              �?      �?        ۶m۶m�?�$I�$I�?              �?C��6�S�?�}�K�`�?�q�q�?�q�q�?      �?        I�$I�$�?۶m۶m�?      �?        F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?        <<<<<<�?�?      �?      �?۶m۶m�?�$I�$I�?�?�?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?�������?333333�?      �?              �?      �?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�;hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������       V                    �?��l�Qf�?�           8�@                                    @�������?�            �p@                                 �;@BӀN��?[            �b@                                  �:@Xny��?$            �N@                                 �7@ �h�7W�?!            �J@       ������������������������       �                     B@                                    �?@�0�!��?
             1@        ������������������������       �                     "@        	       
                   �+@      �?              @        ������������������������       �                     @        ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?                                  �/@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                   �?�E�����?7            �V@                                  �?`����֜?*            �Q@                                  �H@P���Q�?             4@       ������������������������       �        	             (@                                   J@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     I@        ������������������������       �                     4@               O                 03�7@\X��t�?I            �\@              H                 ��.@J`mL�#�?;            @X@              5                 pF @v�(��O�?-            �R@              &                    �?�GN�z�?             F@              %                    �?PN��T'�?             ;@                                �|Y8@HP�s��?             9@        ������������������������       �                     @        !       $                 ���@�C��2(�?             6@        "       #                 �Y�@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             1@        ������������������������       �                      @        '       (                  s@ҳ�wY;�?             1@        ������������������������       �                      @        )       .                 �&B@���Q��?
             .@        *       +                    4@      �?             @        ������������������������       �                      @        ,       -                 �|Y:@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        /       0                 P�@�q�q�?             "@        ������������������������       �                      @        1       4                    �?և���X�?             @       2       3                   �9@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        6       ;                   �1@¦	^_�?             ?@        7       8                    �?      �?              @        ������������������������       �                     @        9       :                    @���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        <       A                 �|�=@�LQ�1	�?             7@       =       >                 �?�-@��S�ۿ?	             .@       ������������������������       �                     &@        ?       @                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        B       C                    �?      �?              @        ������������������������       �                     @        D       E                  SE"@�q�q�?             @        ������������������������       �                     �?        F       G                   &@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       J                    �?�C��2(�?             6@        ������������������������       �                     (@        K       N                    �?z�G�z�?             $@       L       M                 �|�;@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        P       S                    @�����H�?             2@        Q       R                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        T       U                    @      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        W       ^                    *@R�����?           �{@        X       Y                 �Q��?�X����?             6@        ������������������������       �                     @        Z       [                    �?b�2�tk�?
             2@        ������������������������       �                     @        \       ]                   �;@��S���?	             .@        ������������������������       �                      @        ������������������������       �                     @        _       �                    �?�����?           pz@        `       e                   �7@��s����?1             U@        a       d                 ���A@      �?              @       b       c                    5@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        f       �                 �̾w@$�Z����?,             S@       g       �                    �?�r����?+            �R@       h       i                   @@؇���X�?(            �Q@        ������������������������       �                     6@        j       w                 �|Y=@�q�q�?             H@        k       r                     @�eP*L��?	             &@       l       q                     �?�q�q�?             @       m       p                    �?���Q��?             @       n       o                   �8@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        s       v                    <@���Q��?             @       t       u                 �0@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        x       �                     �?$G$n��?            �B@       y       �                    �?"pc�
�?             6@       z       �                   �H@�<ݚ�?             2@       {       ~                 ��2>@�	j*D�?             *@        |       }                 ���<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               �                    C@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��S�ۿ?             .@       ������������������������       �                     (@        �       �                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                     �?��u2��?�            0u@        �       �                   �>@x��}�?$            �K@        �       �                 �|Y<@p�ݯ��?             3@        ������������������������       �                      @        �       �                   @=@�t����?             1@       �       �                 ��<:@z�G�z�?
             .@        ������������������������       �                     @        �       �                 �|�?@�q�q�?             "@        ������������������������       �                     @        �       �                 `f�;@      �?             @       �       �                   @I@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?r�q��?             B@       �       �                   �E@z�G�z�?             >@       �       �                   �B@ҳ�wY;�?             1@       �       �                 �|�<@d}h���?
             ,@        �       �                 `f�D@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 `f�K@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                     @        �       �                 0�H@@�j;��?�            �q@       �       �                    �?�E�J��?�            �p@       �       �                    �?X����?�            `o@        �       �                 �|Y=@$G$n��?            �B@        ������������������������       �                      @        �       �                 X��A@�#-���?            �A@       �       �                   `3@ףp=
�?             >@       �       �                 ���@ 	��p�?             =@        ������������������������       �                     @        �       �                 ��(@�C��2(�?             6@       ������������������������       �      �?	             0@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @tCo���?�            �j@        �       �                 `f�)@@��8��?              H@        ������������������������       �                     4@        �       �                    ,@h�����?             <@        �       �                   @D@$�q-�?	             *@       ������������������������       �                     $@        �       �                   �F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        �       �                 �|�=@�}#���?o            �d@       �       �                   �;@��GEI_�?R            �^@       �       �                   �:@p`q�q��?2            �S@       �       �                 pf� @��S�ۿ?0            �R@       �       �                   �2@ףp=
�?"             I@        ������������������������       �                     $@        �       �                 �?�@      �?             D@       �       �                 ���@`Jj��?             ?@        �       �                 ���@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     7@        �       �                 @3�@�q�q�?             "@        �       �                   �4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �4@�q�q�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     9@        �       �                 �� @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �|Y=@ qP��B�?             �E@        ������������������������       �                     $@        �       �                 ��) @Pa�	�?            �@@       ������������������������       �                     6@        �       �                 pf� @�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 �?�@��2(&�?             F@        ������������������������       �                     5@        �       �                 @3�@��+7��?             7@        �       �                   �?@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �A@      �?              @       ������������������������       ����Q��?             @        ������������������������       ��q�q�?             @        �       �                    ?@@4և���?
             ,@        �       �                 �̌!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     2@        �       �                     @������?             .@        ������������������������       �                      @        �       �                    �?�	j*D�?             *@       �       �                 �|�>@���Q��?             $@       �       �                    ;@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������}<����?�/���?��9����?\�qA��?ـl@6 �?�7���M�?�}�K�`�?C��6�S�?"5�x+��?��sHM0�?              �?�������?ZZZZZZ�?              �?      �?      �?      �?                      �?      �?      �?              �?�$I�$I�?۶m۶m�?              �?      �?        l�l��?P��O���?�A�A�?�������?�������?ffffff�?              �?      �?      �?      �?                      �?              �?              �?��Moz��?!Y�B�?�'�i�n�?5l7˓��?O贁N�?Y�%�X�?]t�E�?�袋.��?h/�����?&���^B�?{�G�z�?q=
ףp�?              �?F]t�E�?]t�E�?�������?333333�?              �?      �?                      �?      �?        �������?�������?              �?�������?333333�?      �?      �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?333333�?�������?      �?                      �?              �?��Zk���?�RJ)���?      �?      �?              �?�������?333333�?              �?      �?        ��Moz��?Y�B��?�������?�?      �?              �?      �?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?F]t�E�?]t�E�?              �?�������?�������?      �?      �?      �?                      �?              �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?      �?      �?                      �?�'�R0�?9a��>��?]t�E]�?�E]t��?              �?9��8���?�8��8��?              �?�������?�?              �?      �?        4F���?��/�	�?z��y���?�a�a�?      �?      �?      �?      �?      �?                      �?              �?�5��P^�?l(�����?�������?�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?�������?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?333333�?�������?      �?      �?      �?                      �?      �?              �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?к����?���L�?/�袋.�?F]t�E�?9��8���?�q�q�?vb'vb'�?;�;��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?                      �?      �?              �?        �������?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?5�M��?Y����?pX���o�?A��)A�?^Cy�5�?Cy�5��?              �?�������?�������?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?�������?333333�?              �?      �?              �?                      �?�������?UUUUUU�?�������?�������?�������?�������?I�$I�$�?۶m۶m�?333333�?�������?              �?      �?        �q�q�?�q�q�?      �?                      �?              �?      �?              �?        w�'�K�?H���@��?�-���?��~���?�_FA@s�?���e�?к����?���L�?              �?�A�A�?_�_�?�������?�������?������?�{a���?      �?        ]t�E�?F]t�E�?      �?      �?      �?                      �?      �?        
�N]���?�_���?UUUUUU�?UUUUUU�?      �?        �m۶m��?�$I�$I�?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        Y1P�M�?4u~�!��?�d����?;ڼOqɰ?T:�g *�?^-n����?�������?�?�������?�������?      �?              �?      �?���{��?�B!��?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?              �?      �?      �?                      �?��}A�?�}A_З?      �?        |���?|���?      �?        ]t�E�?F]t�E�?              �?      �?        ��.���?t�E]t�?      �?        zӛ����?Y�B��?�q�q�?r�q��?              �?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        wwwwww�?�?      �?        vb'vb'�?;�;��?333333�?�������?۶m۶m�?�$I�$I�?              �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ� �thG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                 `fK@���*1�?�           8�@              e                 `f�$@J��u�?}           ��@                                    �?h�3A_'�?�            pp@                                   �?��Sݭg�?            �C@                                �|�9@�t����?             1@        ������������������������       �                     @               
                 ���@8�Z$���?	             *@               	                 �Y�@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@                                   �?���|���?             6@                                  �?���Q��?             4@                               P�@b�2�tk�?             2@                                   4@"pc�
�?             &@        ������������������������       �                     �?                                ���@ףp=
�?             $@        ������������������������       �                     @                                  �A@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   3@����X�?             @        ������������������������       �                     �?                                ��� @r�q��?             @        ������������������������       �                     @                                   :@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                  �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        !       4                    �?@4և���?�             l@        "       1                 ��i @�θ�?             :@       #       *                 �|Y=@�q�q�?             8@        $       %                    5@���Q��?             $@        ������������������������       �                     @        &       '                 ���@z�G�z�?             @        ������������������������       �                      @        (       )                   @@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        +       0                 �|�=@@4և���?             ,@       ,       -                 ���@      �?              @        ������������������������       �                     @        .       /                   @@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        2       3                 Ь:!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        5       D                   �<@ ���v��?y            �h@        6       7                    �? qP��B�?3            �U@        ������������������������       �                      @        8       C                   �4@�Ń��̧?2             U@        9       :                 �?�@�X�<ݺ?             B@        ������������������������       �        
             0@        ;       <                   �1@ףp=
�?             4@        ������������������������       �                     @        =       >                   �2@�r����?             .@        ������������������������       �                     �?        ?       @                   �3@@4և���?             ,@        ������������������������       �                      @        A       B                 @3�@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     H@        E       b                 ���"@@4և���?F             \@       F       G                  s�@�X�<ݺ?D             [@        ������������������������       �                     G@        H       [                 @3�@��a�n`�?*             O@       I       X                 �?�@��hJ,�?             A@       J       M                 �|Y=@ףp=
�?             >@        K       L                   @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        N       O                    �?@4և���?             <@        ������������������������       �                     $@        P       W                   @@@�����H�?             2@       Q       V                   �@8�Z$���?	             *@        R       U                 �&B@�q�q�?             @       S       T                 �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        Y       Z                   �A@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        \       a                 �|�>@h�����?             <@       ]       ^                 ��) @��S�ۿ?
             .@       ������������������������       �                     *@        _       `                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        c       d                 �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        f       �                 `f�:@�M�Ta5�?�            u@       g       �                    :@ҲW��?�            �l@       h       �                    �?�-����?�             k@       i       t                   �;@ (�^G�?^            �a@        j       o                    �?؇���X�?            �A@        k       l                    �?���Q��?             @        ������������������������       �                      @        m       n                     @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        p       s                    4@��S�ۿ?             >@        q       r                   �2@r�q��?             (@       ������������������������       �                     "@        ������������������������       ��q�q�?             @        ������������������������       �                     2@        u       �                 pff/@�q�q�?G             [@       v                           �?:���W�?'            �M@        w       x                 `f�)@�LQ�1	�?             7@        ������������������������       �                      @        y       z                   �B@z�G�z�?
             .@       ������������������������       �                      @        {       |                    D@և���X�?             @        ������������������������       �                      @        }       ~                    ,@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?������?             B@        ������������������������       �                     @        �       �                   �*@XB���?             =@       �       �                 `f�)@�}�+r��?             3@       ������������������������       �                     "@        �       �                   �C@ףp=
�?             $@        ������������������������       �                     @        �       �                   �G@r�q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?�`���?             �H@        �       �                     @�8��8��?             8@       ������������������������       �                     (@        �       �                 03�1@r�q��?             (@       ������������������������       �                     "@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|�=@HP�s��?             9@        �       �                  �v6@�<ݚ�?             "@       ������������������������       �                     @        �       �                    �?      �?             @       �       �                 03�7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                     @z�7�Z�?,            @R@        �       �                    �?ףp=
�?             4@       ������������������������       �                     ,@        �       �                   `6@�q�q�?             @        ������������������������       �                      @        �       �                   �3@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?��k��?             �J@       �       �                    �?��S���?             >@        �       �                 `�@1@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                   �*@և���X�?             5@        ������������������������       �                     @        �       �                 `f7@X�Cc�?             ,@       �       �                 ��/@      �?             $@        ������������������������       �                     @        �       �                    �?����X�?             @       �       �                   �3@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|Y?@�LQ�1	�?             7@       �       �                    �?�t����?
             1@       �       �                    @r�q��?             (@        ������������������������       �                     �?        �       �                 `f2@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �J@z�G�z�?	             .@       �       �                    �?؇���X�?             ,@       �       �                 �|�?@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �3@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �J@���vq�?D            �Z@       �       �                 ��i=@6n�
$)�?<            �W@        �       �                    �?�����?             5@        �       �                 03�;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             1@        �       �                     @�!�,�E�?0            @R@       �       �                    �?��e�B��?#            �I@       �       �                    �?��
ц��?            �C@        ������������������������       �                      @        �       �                   �H@�4�����?             ?@       �       �                 �|Y<@�c�Α�?             =@        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     �?z�G�z�?             9@       �       �                 �|Y>@�q�q�?             8@        �       �                  Y>@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                   @C@؇���X�?	             ,@        ������������������������       �                      @        �       �                 �TA@@�q�q�?             @        ������������������������       �                     �?        �       �                  x#J@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?r�q��?
             (@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                 pV�C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @��2(&�?             6@        �       �                    �?և���X�?             @        ������������������������       �                     @        �       �                 ��T?@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             .@        ������������������������       �                     (@        �                         �N@���"͏�?F            �[@       �       �                    �?�<ݚ�?D             [@       �       �                    �?����e��?*            �P@       ������������������������       �        $             K@        �       �                     @�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?               	                   �?��6���?             E@                                �8@�	j*D�?
             *@                                 �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                              xCQ@      �?              @                                 I@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        
                      03�M@J�8���?             =@                                   @      �?              @        ������������������������       �                      @                                 >@r�q��?             @                                ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �?؇���X�?             5@                                �?�}�+r��?
             3@        ������������������������       �                     �?                                 �?�X�<ݺ?	             2@                                H@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������`l����??'��d�?:m���?�%�X��?��S��?���'���?�i�i�?�|˷|��?�?<<<<<<�?              �?;�;��?;�;��?      �?      �?              �?      �?                      �?F]t�E�?]t�E]�?�������?333333�?9��8���?�8��8��?F]t�E�?/�袋.�?      �?        �������?�������?              �?�������?�������?              �?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?                      �?n۶m۶�?�$I�$I�?ى�؉��?�؉�؉�?UUUUUU�?�������?333333�?�������?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?n۶m۶�?�$I�$I�?      �?      �?      �?              �?      �?      �?      �?      �?              �?              �?      �?              �?      �?        �y;Cb�?1ogH�۩?��}A�?�}A_З?      �?        ��<��<�?�a�a�?��8��8�?�q�q�?      �?        �������?�������?      �?        �������?�?              �?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        n۶m۶�?�$I�$I�?��8��8�?�q�q�?      �?        �s�9��?�c�1Ƹ?KKKKKK�?�������?�������?�������?      �?      �?              �?      �?        n۶m۶�?�$I�$I�?      �?        �q�q�?�q�q�?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?              �?              �?      �?      �?        UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?�������?�?      �?              �?      �?      �?                      �?      �?              �?      �?              �?      �?        �l!�-��?�&�פ��?�Cł��?��xu�2�?�Kh/��?�Kh/���?������?9 2ܫ`�?۶m۶m�?�$I�$I�?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?_[4��?A�Iݗ��?Y�B��?��Moz��?              �?�������?�������?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?        �q�q�?�q�q�?      �?        GX�i���?�{a���?�5��P�?(�����?      �?        �������?�������?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        ����S�?և���X�?UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        q=
ףp�?{�G�z�?9��8���?�q�q�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �lٲe��?�I�&M��?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        "5�x+��?oe�Cj��?�?�������?9��8���?�q�q�?      �?                      �?۶m۶m�?�$I�$I�?              �?%I�$I��?�m۶m��?      �?      �?      �?        �$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?      �?        d!Y�B�?Nozӛ��?�?<<<<<<�?UUUUUU�?�������?      �?        F]t�E�?]t�E�?              �?      �?                      �?      �?        �������?�������?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?      �?      �?              �?      �?      �?              �?      �?              �?        ��}�	�?�����?�+����?ڨ�l�w�?=��<���?�a�a�?      �?      �?              �?      �?              �?        �&M�4i�?ٲe˖-�?�������?�������?�;�;�?�؉�؉�?              �?���Zk��?��RJ)��?5�rO#,�?�{a���?      �?      �?              �?      �?      �?      �?                      �?�������?�������?UUUUUU�?�������?ffffff�?333333�?              �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?                      �?UUUUUU�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?��.���?t�E]t�?�$I�$I�?۶m۶m�?      �?              �?      �?      �?                      �?      �?              �?        *�Y7�"�?v�)�Y7�?�q�q�?9��8���?|���?�>����?              �?UUUUUU�?UUUUUU�?              �?      �?        b�a��?=��<���?;�;��?vb'vb'�?333333�?�������?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�rO#,��?|a���?      �?      �?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?�5��P�?(�����?      �?        ��8��8�?�q�q�?�������?�?      �?                      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��1hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       p                     @�,�٧��?�           8�@               _                    �?0Z� ���?�            ps@              D                     �?Pr=x)��?�            �l@               #                  x#J@j���� �?I            �]@               "                   �M@�0u��A�?$             N@                                  �?z�):���?             I@               
                    �?d}h���?             ,@               	                   �H@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                �|�<@�q�q�?             B@                                `f�D@����X�?             @       ������������������������       �                     @        ������������������������       �                      @               !                 �TA@@>���Rp�?             =@                               ��I/@     ��?             0@        ������������������������       �                     @                                   �?��
ц��?
             *@                                 �>@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                   �>@X�<ݚ�?             "@                               `f�<@      �?              @                               03k:@      �?             @        ������������������������       �                     �?                                   H@���Q��?             @        ������������������������       �                      @                                  �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     $@        $       -                   �4@$gv&��?%            �M@        %       *                    �?      �?              @        &       '                 �U�X@���Q��?             @        ������������������������       �                     �?        (       )                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        +       ,                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        .       A                  �k@>a�����?            �I@       /       6                    B@�LQ�1	�?             G@       0       5                   �9@h�����?             <@        1       4                 0wKT@؇���X�?             @        2       3                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        7       >                 ��Q@�E��ӭ�?             2@       8       9                    C@���Q��?             $@        ������������������������       �                      @        :       ;                    �?      �?              @        ������������������������       �                      @        <       =                 ��DM@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ?       @                   @G@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        B       C                 X�,@@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        E       R                    �?�>4ևF�?L             \@        F       M                   �;@Du9iH��?            �E@        G       H                    �?����X�?             @        ������������������������       �                      @        I       J                   �5@���Q��?             @        ������������������������       �                      @        K       L                   �'@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        N       O                   �E@������?             B@       ������������������������       �                     ;@        P       Q                    5@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        S       T                   �)@�nkK�?2            @Q@        ������������������������       �                     ;@        U       ^                   @A@@4և���?             E@       V       ]                 ��,@ȵHPS!�?             :@        W       X                 �|�<@      �?	             (@       ������������������������       �                     @        Y       Z                 �|�=@      �?             @        ������������������������       �                      @        [       \                    @@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �        	             ,@        ������������������������       �                     0@        `       e                    �?��Q���?4             T@       a       d                    @`Ql�R�?             �G@        b       c                     �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �F@        f       m                 0�X@���|���?            �@@       g       h                    +@j���� �?             1@        ������������������������       �                     "@        i       j                 ��UO@      �?              @       ������������������������       �                     @        k       l                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        n       o                   �4@      �?             0@        ������������������������       �                      @        ������������������������       �                     ,@        q       �                  �#@&S��:�?�             y@       r       �                    �?@�0�!��?�            �o@        s       �                 pF @�zv�X�?             F@       t       u                    �?������?             A@       ������������������������       �        
             0@        v       �                    ;@X�<ݚ�?	             2@       w       �                    �?�θ�?             *@       x       }                   �6@      �?             (@       y       |                   �2@      �?              @        z       {                 P��@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ~                          �8@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �3@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?�S	���?�            `j@        �       �                    �?��E�B��?            �G@       �       �                    �?�����H�?            �F@        �       �                   �6@���}<S�?             7@        ������������������������       �                      @        ������������������������       �                     5@        �       �                 �|Y=@��2(&�?             6@        �       �                  ��@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                  s�@�KM�]�?             3@        ������������������������       �                     @        ������������������������       �؇���X�?	             ,@        �       �                 ��}@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|�=@��p\�?e            �d@       �       �                 �?$@ \sF��?F            @\@        �       �                 ��@$�q-�?            �C@       �       �                    7@�g�y��?             ?@       ������������������������       �        
             0@        �       �                 ���@��S�ۿ?             .@        �       �                   `@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 �|�;@      �?              @       ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                   �2@�?�|�?/            �R@        �       �                 ��Y @r�q��?             (@        �       �                    1@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �        )             O@        �       �                   �"@L紂P�?            �I@       �       �                 �?�@dP-���?            �G@       ������������������������       �                     <@        �       �                 @3�@���y4F�?             3@        �       �                   �?@      �?              @        ������������������������       �                     �?        �       �                   �A@և���X�?             @       ������������������������       ��q�q�?             @        ������������������������       �      �?             @        ������������������������       �                     &@        �       �                   �?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                  ��8@20J�Ws�?Y             b@       �       �                    �?�~8�e�?>            �Y@        �       �                    �?d,���O�?            �I@        �       �                    �?؇���X�?             <@       �       �                 pF�-@H%u��?             9@        �       �                    >@      �?             (@       �       �                 P��+@"pc�
�?             &@        ������������������������       �                     @        �       �                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @�û��|�?             7@        ������������������������       �                     @        �       �                 �|�<@      �?             2@       �       �                    �?�z�G��?             $@       �       �                    4@      �?              @       �       �                 `F�+@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �C@      �?              @       �       �                   �>@؇���X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    $@x�K��?!            �I@        ������������������������       �                     $@        �       �                 ��-@���?            �D@        �       �                    �?��S�ۿ?
             .@        �       �                    3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                 ��.@$��m��?             :@        ������������������������       �                     @        �       �                 03�6@�GN�z�?             6@       �       �                    �?r�q��?             2@       ������������������������       �        
             (@        �       �                 8#"2@      �?             @        �       �                    >@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?X�EQ]N�?            �E@        ������������������������       �                     @        �       �                    �?4?,R��?             B@        ������������������������       �                      @        �       �                    �?�>4և��?             <@       �       �                 ��p@@�KM�]�?             3@        �       �                     @�<ݚ�?             "@        �       �                    @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    @�q�q�?             "@       �       �                    @      �?              @        �       �                     @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������&��jq�?:�g *�?AW o��?_��oH��?�bAs�X�?�:}�N�?ZZZZZZ�?�������?�������?�������?H�z�G�?q=
ףp�?۶m۶m�?I�$I�$�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?�$I�$I�?�m۶m��?              �?      �?        �i��F�?GX�i���?      �?      �?      �?        �؉�؉�?�;�;�?      �?      �?      �?                      �?�q�q�?r�q��?      �?      �?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?              �?        ��/���?[4��}�?      �?      �?333333�?�������?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �?�������?Y�B��?��Moz��?�$I�$I�?�m۶m��?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?r�q��?�q�q�?�������?333333�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?�������?333333�?      �?                      �?n۶m۶�?%I�$I��?w�qGܱ?qG�w��?�$I�$I�?�m۶m��?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?              �?�q�q�?�q�q�?              �?      �?        �Mozӛ�?d!Y�B�?      �?        n۶m۶�?�$I�$I�?��N��N�?�؉�؉�?      �?      �?      �?              �?      �?              �?      �?      �?      �?              �?      �?      �?              �?        �������?333333�?W�+�ɕ?}g���Q�?      �?      �?      �?                      �?              �?]t�E]�?F]t�E�?ZZZZZZ�?�������?              �?      �?      �?      �?              �?      �?              �?      �?              �?      �?              �?      �?        \���(\�?H�z�G�?ZZZZZZ�?�������?�袋.��?��.���?�?xxxxxx�?              �?�q�q�?r�q��?�؉�؉�?ى�؉��?      �?      �?      �?      �?�������?�������?              �?      �?                      �?      �?      �?      �?                      �?              �?      �?        �������?�������?              �?      �?        �ƴ	(E�?1�Y��ֵ?�l�w6��?AL� &W�?�q�q�?�q�q�?ӛ���7�?d!Y�B�?              �?      �?        ��.���?t�E]t�?UUUUUU�?UUUUUU�?      �?                      �?�k(���?(�����?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?�]�ڕ��?��+Q��?[X驅��?Vzja���?�؉�؉�?;�;��?��{���?�B!��?      �?        �������?�?      �?      �?      �?                      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?*�Y7�"�?к����?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        �������?�������?�����F�?W�+�ɵ?      �?        6��P^C�?(������?      �?      �?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?              �?      �?        z�!���?�Ő��?�������?222222�?PPPPPP�?�������?�$I�$I�?۶m۶m�?���Q��?)\���(�?      �?      �?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ��,d!�?8��Moz�?              �?      �?      �?ffffff�?333333�?      �?      �?      �?      �?              �?      �?              �?              �?              �?      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ssssss�?�?              �?28��1�?8��18�?�������?�?UUUUUU�?UUUUUU�?              �?      �?              �?        �N��N��?vb'vb'�?              �?�袋.��?]t�E�?�������?UUUUUU�?      �?              �?      �?      �?      �?              �?      �?              �?              �?      �?              �?      �?        w�qG�?qG�wĽ?      �?        �8��8��?r�q��?      �?        �$I�$I�?�m۶m��?�k(���?(�����?9��8���?�q�q�?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?      �?      �?�������?333333�?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�JIhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       H                     �?���*1�?�           8�@                                   �?2p�ZAJ�?e            �c@                                   �?�b��-8�?(            �O@        ������������������������       �                     @@                                p"�X@`՟�G��?             ?@                                  �?�q�����?             9@                                xCH@���Q��?             4@              	                 `f&;@���!pc�?             &@        ������������������������       �                     �?        
                        �|�=@z�G�z�?             $@                                ��2>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   C@      �?              @        ������������������������       �                     @                                  �H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@                                ��UO@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?r�q��?             @        ������������������������       �                     @                                  �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               9                 ��gS@�q�q�?=             X@              8                 03�M@TV����?&            �M@                                  �?䯦s#�?#            �J@        ������������������������       �                     $@                7                    K@v ��?            �E@       !       "                 �̌*@�e����?            �C@        ������������������������       �                     @        #       $                    7@*O���?             B@        ������������������������       �                      @        %       &                   �<@�!���?             A@        ������������������������       �                     @        '       0                   `@@�5��?             ;@        (       )                 �|Y=@������?             1@        ������������������������       �                     @        *       /                 `fF<@@4և���?             ,@       +       .                   @G@z�G�z�?             @        ,       -                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        1       2                  x#J@�z�G��?             $@       ������������������������       �                     @        3       6                   �C@      �?             @       4       5                    A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        :       =                    �?�MI8d�?            �B@        ;       <                   @C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        >       E                  �k@�C��2(�?            �@@       ?       @                    �?(;L]n�?             >@       ������������������������       �                     8@        A       D                    F@r�q��?             @       B       C                    5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        F       G                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        I       �                    �?�q�q�?W           @�@        J       W                    �?���#��?i            �d@        K       N                   �-@$G$n��?            �B@        L       M                 `�@1@      �?             @        ������������������������       �                     @        ������������������������       �                     @        O       R                 ���@`Jj��?             ?@        P       Q                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       T                    �?XB���?             =@       ������������������������       �                     ;@        U       V                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        X       o                  �#@B@��S��?M             `@        Y       j                   �7@���Q��?            �A@       Z       c                   �5@և���X�?             5@       [       \                 ���@���|���?             &@        ������������������������       �                     @        ]       `                   �2@և���X�?             @        ^       _                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        a       b                    4@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        d       g                   �6@      �?             $@       e       f                 �̜!@      �?              @       ������������������������       �                     @        ������������������������       �                     @        h       i                 @3�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        k       l                 �|Y>@؇���X�?             ,@       ������������������������       �                      @        m       n                    A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        p       �                 03�>@z�J�?:            �W@       q       �                    @h/��y��?,            @S@       r       �                     @�d�����?+             S@       s       �                    :@��2(&�?             F@       t       �                   �J@�n`���?             ?@       u       v                   �'@r�q��?             >@        ������������������������       �                     (@        w       �                    �?�E��ӭ�?             2@       x       }                   �7@      �?	             $@       y       z                   �<@�q�q�?             @        ������������������������       �                     @        {       |                   �A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ~                          @B@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    @     ��?             @@        ������������������������       �                     @        �       �                 03�1@|��?���?             ;@       �       �                    �?������?             1@       �       �                 ��&@@4և���?             ,@        �       �                 �[$@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        �       �                     @ҳ�wY;�?             1@        ������������������������       �                     @        �       �                    @�8��8��?	             (@       ������������������������       �                      @        �       �                   @C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@��y�S��?�             x@        �       �                 �|Y=@,�d�vK�?X            �a@        �       �                 ��@(N:!���?+            �Q@       �       �                   �<@"pc�
�?            �@@       �       �                   �3@��� ��?             ?@        ������������������������       �                      @        �       �                    �?�㙢�c�?             7@        �       �                   �6@����X�?             @        �       �                 ��y@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    7@      �?
             0@       ������������������������       �                     "@        �       �                 ���@����X�?             @        �       �                 �&b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?@-�_ .�?            �B@       �       �                   �<@ >�֕�?            �A@       ������������������������       �                    �@@        ������������������������       �                      @        ������������������������       �                      @        �       �                     @ �q�q�?-             R@        ������������������������       �                     �?        �       �                    �?0z�(>��?,            �Q@       �       �                 ���@������?             B@        �       �                 ���@$�q-�?             *@       ������������������������       �                     "@        �       �                 �|�=@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     7@        �       �                 �&B@ >�֕�?            �A@        ������������������������       �                     6@        �       �                    ?@8�Z$���?
             *@       ������������������������       �                     @        �       �                   �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �4@yٯ���?�            �n@        �       �                 0S5 @�d�K���?+            �P@        �       �                 @3�@d}h���?             ,@        ������������������������       ��q�q�?             @        �       �                   �3@"pc�
�?             &@       �       �                    1@ףp=
�?             $@        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���$@�q����?$            �J@        �       �                 �-!@�X�<ݺ?             2@        �       �                ��k"@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                     @և���X�?            �A@        �       �                    �?����X�?             @        �       �                    &@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 03�0@X�Cc�?             <@        ������������������������       �                     "@        �       �                 `f68@�}�+r��?             3@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                     @(+���?k             f@        �       �                 �|�=@`׀�:M�?)            �R@        �       �                    �?@4և���?
             ,@       �       �                 ��,@$�q-�?	             *@       �       �                 �|�<@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     N@        �       �                 @3�@=�Ѝ;�?B            �Y@        �       �                    >@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �                          �?<����?>            �W@       �       �                 ��q1@�:�^���?;            �V@       �       �                 �|�=@ �q�q�?/             R@       �       �                 ��-@`Ql�R�?            �G@       ������������������������       �                     C@        �       �                 ��.@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��)"@HP�s��?             9@       ������������������������       �                     0@        �       �                    �?�<ݚ�?             "@       �       �                   �?@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�E��ӭ�?             2@        �       �                 �|�;@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �T)D@؇���X�?
             ,@       ������������������������       �                     $@                                  ;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������`l����??'��d�?Eg@(��?]z��k#�?QEQE�?�u]�u]�?              �?�1�c��?�s�9��?���Q��?�p=
ף�?�������?333333�?F]t�E�?t�E]t�?              �?�������?�������?      �?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?                      �?�������?�������?      �?                      �?�������?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?u_[4�?E�pR���?�V�9�&�?�����?              �?qG�w��?G�w��?�A�A�?�-��-��?      �?        �q�q�?�q�q�?      �?        �������?�������?              �?/�����?h/�����?�?xxxxxx�?      �?        �$I�$I�?n۶m۶�?�������?�������?      �?      �?              �?      �?                      �?              �?ffffff�?333333�?      �?              �?      �?      �?      �?              �?      �?                      �?      �?              �?        L�Ϻ��?��L���?      �?      �?              �?      �?        F]t�E�?]t�E�?�?�������?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?%�����?~�!��?���L�?к����?      �?      �?      �?                      �?�B!��?���{��?      �?      �?              �?      �?        �{a���?GX�i���?              �?      �?      �?              �?      �?        sƜ1g��?Ɯ1g��?333333�?�������?۶m۶m�?�$I�$I�?F]t�E�?]t�E]�?              �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?              �?      �?              �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �w6�;�?��
br�?V~B����?���15��?y�5���?Cy�5��?t�E]t�?��.���?�c�1��?�9�s��?UUUUUU�?�������?              �?r�q��?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?                      �?      �?                      �?      �?      �?              �?{	�%���?	�%����?�?xxxxxx�?�$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?      �?              �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �l.j��?�LF�W>�?��9�h��?�z2~�Գ?|�W|�W�?�A�A�?/�袋.�?F]t�E�?�{����?�B!��?      �?        �7��Mo�?d!Y�B�?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?              �?      �?      �?        �m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?                      �?S�n0E�?к����?��+��+�?�A�A�?      �?                      �?      �?        �������?UUUUUU�?      �?        �ԓ�ۥ�?H���@��?�q�q�?�q�q�?�؉�؉�?;�;��?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        ��+��+�?�A�A�?      �?        ;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?        �u�y��?��).��?�rv��?����?۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?F]t�E�?/�袋.�?�������?�������?�������?�������?              �?      �?        �Cj��V�?�x+�R�?��8��8�?�q�q�?�������?UUUUUU�?              �?      �?              �?        �$I�$I�?۶m۶m�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?%I�$I��?�m۶m��?              �?�5��P�?(�����?�������?�������?      �?                      �?      �?        �?�x�?�^o�?�?��L��?к����?n۶m۶�?�$I�$I�?�؉�؉�?;�;��?۶m۶m�?�$I�$I�?      �?                      �?      �?              �?              �?        ������?R�yY�'�?      �?      �?      �?                      �?���%N�?�X�0Ҏ�?}�'}�'�?l�l��?�������?UUUUUU�?}g���Q�?W�+�ɕ?      �?        �q�q�?�q�q�?              �?      �?        q=
ףp�?{�G�z�?      �?        9��8���?�q�q�?333333�?�������?              �?      �?              �?        �q�q�?r�q��?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��NhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       \                 `f�%@���%&�?�           8�@               )                    �?�DgdK+�?�            r@                                `��!@�u���?&            �N@                                  �?���X�K�?            �F@                                   �?R���Q�?             4@        ������������������������       �                     �?               
                    �?�S����?             3@              	                 ���@�����H�?
             2@        ������������������������       �                      @        ������������������������       �        	             0@        ������������������������       �                     �?                                �&B@���Q��?             9@                                   8@�q�q�?             "@                               pf�@���Q��?             @        ������������������������       �                      @                                   4@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                   5@      �?             0@        ������������������������       �                     @                                ��� @���|���?             &@                               P�@      �?              @        ������������������������       �                      @                                  �9@�q�q�?             @        ������������������������       �                     @                                @3�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                    3@     ��?             0@        ������������������������       �                     �?        !       (                    �?������?             .@       "       #                 03S$@�	j*D�?
             *@        ������������������������       �                     @        $       '                   �J@�q�q�?             @       %       &                     @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        *       /                     @l�b�G��?�            �l@        +       ,                     �? �q�q�?             8@        ������������������������       �                     @        -       .                    5@P���Q�?             4@        ������������������������       �      �?             @        ������������������������       �                     0@        0       C                    �?����p�?�            �i@        1       <                  ��@      �?#             L@       2       ;                    �?�IєX�?             A@       3       :                    �?�����?             5@       4       5                 �|=@ףp=
�?             4@        ������������������������       �                     @        6       9                 �|�=@8�Z$���?
             *@       7       8                 ���@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        =       >                 �|Y=@�GN�z�?             6@        ������������������������       �                     @        ?       B                 P�J@�KM�]�?             3@       @       A                 X�I@؇���X�?	             ,@       ������������������������       �r�q��?             (@        ������������������������       �                      @        ������������������������       �                     @        D       E                   �:@@-�_ .�?a            �b@        ������������������������       �        (             P@        F       S                 ��) @�����?9             U@       G       H                   �>@hA� �?0            �Q@        ������������������������       �                     @@        I       J                 �&B@�˹�m��?             C@        ������������������������       �                     4@        K       L                   �@r�q��?             2@        ������������������������       �                     �?        M       N                   �?@�t����?             1@        ������������������������       �                     �?        O       R                 @3�@      �?             0@       P       Q                   @C@�����H�?             "@       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        T       U                 ��y @X�Cc�?	             ,@        ������������������������       �                     @        V       [                 ���!@"pc�
�?             &@       W       X                 pf!@����X�?             @        ������������������������       �                     �?        Y       Z                 �|Y<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ]       �                    �?F7T:`��?           `z@        ^       q                     @�����?�             i@       _       f                   �E@����Q8�?X            �a@       `       a                    �?�]���?J            �\@        ������������������������       �                    �B@        b       c                    :@ ���J��?2            �S@        ������������������������       �                     D@        d       e                   �;@�}�+r��?             C@        ������������������������       �                      @        ������������������������       �                     B@        g       p                    �?�<ݚ�?             ;@       h       i                   @F@�q�q�?	             2@        ������������������������       �                     @        j       o                     �?z�G�z�?             .@       k       n                 ��A@d}h���?             ,@        l       m                   �H@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        r       �                 ��Y7@��o	��?(             M@       s       t                 @�+@����X�?            �A@        ������������������������       �                     @        u       �                    �?�q�q�?             >@       v       {                 �?�-@�d�����?             3@        w       x                   �-@�q�q�?             @        ������������������������       �                      @        y       z                   �0@      �?             @        ������������������������       �                      @        ������������������������       �                      @        |       }                    �?$�q-�?	             *@       ������������������������       �                      @        ~       �                    @z�G�z�?             @              �                 �|Y=@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�eP*L��?
             &@       �       �                 �|�<@X�<ݚ�?	             "@       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                    @      �?             @        �       �                 @3�2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @       �       �                 �|Y>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                  ��8@���}<S�?             7@        �       �                 �|�=@      �?             @       �       �                 ���7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�}�+r��?             3@        ������������������������       �                     @        �       �                    @      �?
             0@       ������������������������       �                     ,@        �       �                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                  x#J@"��$�?�            �k@       �       �                    #@�4���L�?l            �e@        �       �                 @3�4@�q�q�?             2@        ������������������������       �                     @        �       �                 ��A>@�eP*L��?             &@       �       �                    @����X�?             @       �       �                     @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @      �?             @       �       �                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?؇���X�?_            @c@       �       �                     �?v���a�?X            @b@        �       �                   �B@ \� ���?!            �H@       �       �                    �?�	j*D�?            �C@       �       �                    �?4�B��?            �B@        �       �                 �|�;@�q�q�?             "@        ������������������������       �                     �?        �       �                  �>@      �?              @       �       �                 X��E@؇���X�?             @       �       �                 �ܵ<@z�G�z�?             @        ������������������������       �                      @        �       �                 ��2>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 `fF:@��X��?             <@        ������������������������       �                     @        �       �                 �TaA@�û��|�?             7@       �       �                  i?@���|���?             6@       �       �                   �J@���Q��?             4@       �       �                 `f�;@�n_Y�K�?             *@       �       �                 �|�?@      �?              @        �       �                 �|�<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   @>@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �                 �|�=@�^'�ë�?7            @X@       �       �                 �&@     ��?             H@        ������������������������       �                     �?        �       �                 �|=@t/*�?            �G@       ������������������������       �                     A@        �       �                    �?�n_Y�K�?             *@       �       �                    �?����X�?             @       �       �                 `fv2@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �+@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �A@@�E�x�?            �H@        �       �                    �?�C��2(�?             &@       �       �                   �@@      �?              @        ������������������������       �                     @        �       �                    1@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     C@        ������������������������       �                      @        �                         @I@� �	��?              I@       �                       �|�>@X��ʑ��?            �E@       �       �                    �?�n_Y�K�?             :@        �       �                   �4@���Q��?             $@        ������������������������       �                     �?        �       �                   �7@�q�q�?             "@        ������������������������       �                     �?        �       �                  �}S@      �?              @        ������������������������       �                     @        �       �                    :@      �?             @       �       �                 0�HU@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �                          �;@      �?
             0@        �       �                   �7@և���X�?             @       �       �                     �?      �?             @       �       �                    '@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@                                �E@�t����?
             1@                              �!fK@�����H�?             "@                              `�iJ@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @              	                  @G@      �?              @        ������������������������       �                      @        
                         �?�q�q�?             @                               �H@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������g *��?�0���M�?�?�0�!�?� =[y�?XG��).�?T\2�h�?�'}�'}�?l�l��?333333�?333333�?              �?^Cy�5�?(������?�q�q�?�q�q�?      �?                      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?F]t�E�?]t�E]�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?wwwwww�?�?vb'vb'�?;�;��?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?              �?        �Gp��?p�}��?�������?UUUUUU�?      �?        ffffff�?�������?      �?      �?      �?        �������?�����Ҳ?      �?      �?�?�?=��<���?�a�a�?�������?�������?      �?        ;�;��?;�;��?9��8���?�q�q�?      �?        333333�?�������?      �?              �?              �?        �袋.��?]t�E�?              �?�k(���?(�����?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?              �?        S�n0E�?к����?      �?        =��<���?�a�a�?���?_�_�?      �?        ��P^Cy�?^Cy�5�?      �?        �������?UUUUUU�?              �?<<<<<<�?�?              �?      �?      �?�q�q�?�q�q�?      �?              �?      �?      �?        %I�$I��?�m۶m��?              �?/�袋.�?F]t�E�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ���X�?,4�Syt�?�(\����?��(\���?��Vج?O�o�z2�?���ϑ?��ʇq�?              �?�A�A�?��-��-�?              �?(�����?�5��P�?      �?                      �?�q�q�?9��8���?UUUUUU�?UUUUUU�?      �?        �������?�������?۶m۶m�?I�$I�$�?      �?      �?              �?      �?                      �?              �?              �?���{�?������?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?y�5���?Cy�5��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ;�;��?�؉�؉�?              �?�������?�������?      �?      �?              �?      �?                      �?]t�E�?t�E]t�?r�q��?�q�q�?�������?�������?      �?              �?      �?      �?      �?              �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?ӛ���7�?d!Y�B�?      �?      �?      �?      �?      �?                      �?      �?        �5��P�?(�����?      �?              �?      �?      �?              �?      �?              �?      �?        �~G����?Nq��$�?kʚ����?S֔5eM�?UUUUUU�?UUUUUU�?              �?t�E]t�?]t�E�?�m۶m��?�$I�$I�?�������?�������?              �?      �?              �?      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?۶m۶m�?�$I�$I�?ٲe˖-�?�4iҤI�?
^N��)�?և���X�?vb'vb'�?;�;��?�Y7�"��?L�Ϻ��?UUUUUU�?UUUUUU�?              �?      �?      �?۶m۶m�?�$I�$I�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?n۶m۶�?%I�$I��?      �?        8��Moz�?��,d!�?]t�E]�?F]t�E�?333333�?�������?ى�؉��?;�;��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?�������?      �?                      �?      �?              �?                      �?      �?              �?        =�L�v��?���Id�?      �?      �?              �?�;����?W�+���?      �?        ى�؉��?;�;��?�$I�$I�?�m۶m��?�������?333333�?              �?      �?                      �?      �?      �?              �?      �?        և���X�?9/���?]t�E�?F]t�E�?      �?      �?      �?              �?      �?      �?      �?      �?              �?              �?              �?        �Q����?)\���(�?��}A�?�}A_�?;�;��?ى�؉��?�������?333333�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?      �?      �?      �?      �?                      �?      �?              �?      �?۶m۶m�?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �������?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?�������?333333�?              �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ2�3hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0Kㅔh2h3h4hph<�h=Kub��������       <                     �?�����?�           8�@                                   �?�`����?h            �d@                                   �?d}h���?,            �Q@                                 �H@����|e�?!             K@                                  �?������?            �B@       ������������������������       �                     9@                                X�,@@�q�q�?	             (@                                Y>@�q�q�?             @        	       
                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                p�9K@��.k���?	             1@       ������������������������       �                     @                                p"W@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @                                 x�E@      �?             0@        ������������������������       �                     �?                                �\@��S�ۿ?
             .@       ������������������������       �                     "@                                   �?r�q��?             @        ������������������������       �                     @                                   C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?               #                    �?�q�q��?<             X@                                ���a@�X�<ݺ?             B@       ������������������������       �                     :@               "                 03c@z�G�z�?             $@                !                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        $       /                   �>@���Q��?%             N@        %       &                 03:@�P�*�?             ?@        ������������������������       �                     @        '       ,                    K@ �o_��?             9@       (       +                   `G@      �?	             0@       )       *                   �F@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        -       .                 `fF<@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        0       1                  x#J@V�a�� �?             =@       ������������������������       �                     1@        2       3                    7@      �?
             (@        ������������������������       �                      @        4       5                   @K@���Q��?	             $@        ������������������������       �                      @        6       7                 �|Y>@      �?              @        ������������������������       �                     �?        8       ;                 03�U@և���X�?             @       9       :                    C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        =       F                    @F�����?S           �@        >       C                    �?     ��?             @@        ?       @                  18@�eP*L��?             &@       ������������������������       �                     @        A       B                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        D       E                 ��yE@���N8�?             5@       ������������������������       �                     4@        ������������������������       �                     �?        G       x                 ���"@P̏����?>           �@        H       I                    /@\�#���?�            �l@        ������������������������       �                     @        J       W                    �?���5��?�            �l@        K       N                    �?d��0u��?             >@        L       M                    �?�r����?	             .@       ������������������������       �                     *@        ������������������������       �                      @        O       V                    �?���Q��?             .@       P       U                   �7@X�Cc�?
             ,@        Q       R                   �6@r�q��?             @       ������������������������       �                     @        S       T                 @3�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        X       i                 �?�@���7�?z            �h@       Y       `                   @4@ ��ʻ��?Y             a@        Z       _                    �? �q�q�?             8@        [       \                 �{@      �?             @        ������������������������       �                      @        ]       ^                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        a       h                    �?����X�?J             \@        b       c                 ���@P���Q�?             4@       ������������������������       �                     (@        d       e                 �|�:@      �?              @        ������������������������       �                      @        f       g                   @@r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �        <             W@        j       k                   �1@X��Oԣ�?!             O@        ������������������������       �                     (@        l       m                   �2@�:pΈ��?             I@        ������������������������       �                      @        n       q                   �4@8��8���?             H@        o       p                 0S @      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        r       w                 @3�@��(\���?             D@        s       t                    >@z�G�z�?             .@        ������������������������       �                     @        u       v                   �A@      �?             (@       ������������������������       �      �?              @        ������������������������       �      �?             @        ������������������������       �                     9@        y       �                    �?Ȅ�<��?�            �q@        z       �                 0C�>@؞�z���?M            @]@       {       �                     @      �?=             V@       |       �                   �E@�NW���?"            �J@       }       ~                   @4@ �q�q�?             H@       ������������������������       �                     ;@               �                   �9@�����?             5@        ������������������������       �                     $@        �       �                   �7@"pc�
�?             &@        �       �                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �G@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��&@��
P��?            �A@        ������������������������       �                     @        �       �                    @     ��?             @@       �       �                   �<@�g�y��?             ?@        �       �                    �?�8��8��?	             (@       ������������������������       �                     $@        �       �                 ��l4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @@���y4F�?             3@       �       �                 �|�=@      �?             0@       �       �                    �?"pc�
�?             &@        �       �                 �|Y=@      �?             @        ������������������������       �                      @        �       �                  S�2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 м[8@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���Q��?             @        �       �                   �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                     @����"�?             =@        ������������������������       �                      @        �       �                 X��@@؇���X�?             5@       ������������������������       �                     &@        �       �                   @C@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                    @lGts��?b            �d@       �       �                    *@�����H�?`            @d@        �       �                 �y.@�	j*D�?             *@        ������������������������       �                     @        �       �                    �?ףp=
�?             $@       ������������������������       �                     @        �       �                 `f68@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     @��7*��?X            �b@       �       �                 �|Y=@P��BNֱ?1            �T@        ������������������������       �                    �@@        �       �                    �? "��u�?             I@        ������������������������       �                     @        �       �                 �|�=@t��ճC�?             F@        ������������������������       �                     �?        �       �                   �@@ �#�Ѵ�?            �E@        ������������������������       �                     ,@        �       �                   @A@ 	��p�?             =@        �       �                    1@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        �       �                    �?`2U0*��?             9@       �       �                   �*@���7�?             6@       �       �                   @D@�8��8��?             (@        ������������������������       �                     @        �       �                   �F@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        �       �                 `�X#@r�q��?'            �P@        �       �                   �8@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?x�}b~|�?#            �L@       �       �                   �3@h�WH��?              K@        ������������������������       �                     .@        �       �                    �?�ݜ�?            �C@        �       �                    �?և���X�?             @       �       �                   �:@���Q��?             @        �       �                 �0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �|�>@      �?             @@       ������������������������       �                     5@        �       �                   @@@�C��2(�?             &@        �       �                 �!B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub������������������?��܍��?�e�@	o�?M�_{��?۶m۶m�?I�$I�$�?	�%����?����K�?к����?��g�`��?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�������?�?      �?        �������?�������?              �?      �?              �?      �?      �?        �?�������?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?�q�q�?��8��8�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?�������?�Zk����?�RJ)���?      �?        �Q����?
ףp=
�?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?��{a�?a���{�?      �?              �?      �?      �?        �������?333333�?              �?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?                      �?4q/;B�?���{��?      �?      �?]t�E�?t�E]t�?              �?�������?UUUUUU�?              �?      �?        �a�a�?��y��y�?              �?      �?        ?���#�?��Gp�?��n���?��D�o-�?              �?�}��?��Gp�?wwwwww�?DDDDDD�?�?�������?              �?      �?        333333�?�������?%I�$I��?�m۶m��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�.�袋�?F]t�E�?�������?�?�������?UUUUUU�?      �?      �?      �?              �?      �?      �?                      �?      �?        n۶m۶�?�$I�$I�?ffffff�?�������?      �?              �?      �?      �?        �������?UUUUUU�?      �?      �?      �?              �?        c�1�c�?�s�9�?      �?        ��Q���?�Q����?              �?�������?�������?      �?      �?UUUUUU�?UUUUUU�?      �?        �������?333333�?�������?�������?      �?              �?      �?      �?      �?      �?      �?      �?        ��şH8�?�2t�n��?^�^��?�P�P�?      �?      �?�x+�R�?萚`���?UUUUUU�?�������?              �?�a�a�?=��<���?              �?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?333333�?      �?                      �?PuPu�?_�_��?      �?              �?      �?��{���?�B!��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        (������?6��P^C�?      �?      �?F]t�E�?/�袋.�?      �?      �?              �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?        �������?333333�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?	�=����?�i��F�?              �?۶m۶m�?�$I�$I�?      �?        ffffff�?333333�?              �?      �?        �<%�S��?�־a�?�q�q�?�q�q�?vb'vb'�?;�;��?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        ]"<)H��?����?��FS���?���ˊ��?      �?        �G�z�?���Q��?      �?        �E]t��?t�E]t�?              �?�/����?�}A_Ч?      �?        ������?�{a���?      �?      �?      �?      �?      �?        ���Q��?{�G�z�?�.�袋�?F]t�E�?UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?              �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?�YLg1�?Lg1��t�?��^B{	�?B{	�%��?      �?        \��[���?�i�i�?۶m۶m�?�$I�$I�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?      �?      �?        ]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJk�ahG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K兔h2h3h4hph<�h=Kub��������       $                    /@	dm#��?�           8�@                                   �?<��¤�?.             Q@                                �&�)@r�q��?             (@        ������������������������       �                     @                                  �,@����X�?             @       ������������������������       �                     @        ������������������������       �                      @                                    @h�����?'             L@        	       
                 �-]@      �?             0@       ������������������������       �                     &@                                   �?z�G�z�?             @                               03�f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                `f7@���Q��?             D@                                   �?r�q��?             2@        ������������������������       �                     @                                   �?z�G�z�?	             .@        ������������������������       �                     �?                                   �?d}h���?             ,@                                  @      �?              @                                  @����X�?             @                                pf�0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                !                 ��T?@���7�?             6@       ������������������������       �        	             (@        "       #                 ��p@@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        %       \                    �?D%���?�           �@        &       [                    @���c�H�?�            �h@       '       <                     @��k=.��?�            �g@       (       -                    �?��p\�?Q            �^@        )       *                   �H@(N:!���?            �A@       ������������������������       �                     8@        +       ,                 83F@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        .       ;                    :@����!p�?;             V@        /       8                   �8@���H��?             E@       0       7                    L@     ��?             @@       1       6                   �9@`Jj��?             ?@        2       3                    5@���Q��?             @        ������������������������       �                      @        4       5                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     :@        ������������������������       �                     �?        9       :                   �E@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        !             G@        =       T                    �?�G\�c�?0            @P@       >       M                 @3�/@θ	j*�?%             J@       ?       F                   �9@0,Tg��?             E@        @       C                  ��@��
ц��?             *@        A       B                   �7@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        D       E                    3@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        G       J                    �?\-��p�?             =@        H       I                 ��%@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        K       L                 ���@$�q-�?             :@        ������������������������       �                      @        ������������������������       �                     8@        N       S                   �4@���Q��?             $@       O       P                 �|�;@      �?              @        ������������������������       �                     @        Q       R                 �|Y>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        U       Z                 �|Y<@�θ�?             *@        V       Y                    �?      �?             @        W       X                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ]       �                     �?���&��?           �{@        ^       �                   �E@�
�G�?9             V@       _       t                    �?П[;U��?#             M@        `       o                   @@@p�ݯ��?             3@       a       n                    �?�eP*L��?
             &@       b       g                 �|�;@      �?	             $@       c       d                    �?z�G�z�?             @       ������������������������       �                     @        e       f                 �nc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        h       m                 �|�=@z�G�z�?             @       i       j                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        k       l                 ��2>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        p       s                 ��Y>@      �?              @        q       r                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        u       �                 �|Y>@�99lMt�?            �C@       v                          �>@�GN�z�?             6@        w       x                 ��<:@���Q��?             $@        ������������������������       �                     @        y       z                   �<@և���X�?             @        ������������������������       �                     @        {       |                 �|Y=@      �?             @        ������������������������       �                     �?        }       ~                 `fF<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �<@�8��8��?             (@        �       �                 `f�D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ��n^@��.k���?             1@       �       �                   �C@�	j*D�?             *@       �       �                   @@@z�G�z�?             $@        �       �                 0��J@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                  �F:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �H@ףp=
�?             >@        �       �                    �?�θ�?	             *@       �       �                   �G@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        �       �                     @p
t�?�            pv@        ������������������������       �        /            @Q@        �       �                   �C@�������?�             r@       �       �                   @C@4Jı@�?�            �o@       �       �                    �?X����?�            `o@        �       �                   �:@     ��?             @@        �       �                    �?�eP*L��?             &@       �       �                 �0@���Q��?             $@       �       �                   �6@�q�q�?             @       �       �                 ��y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�=@؇���X�?             5@       �       �                    �?���!pc�?             &@       �       �                 ��� @�����H�?             "@       �       �                 ��=@z�G�z�?             @        ������������������������       �                     @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?h�j��l�?�            `k@        ������������������������       �                     3@        �       �                 0�H@�Pk�w��?z             i@       �       �                    �?h�a��?v            @h@       �       �                 ���@p�u$v��?n            �f@        ������������������������       �                     4@        �       �                 ���@���`uӽ?c             d@        ������������������������       �                      @        �       �                 �?�@�<� w�?b            �c@        �       �                    ?@P�Lt�<�?,             S@       �       �                 �|�<@@	tbA@�?'            @Q@       ������������������������       �                     H@        �       �                  sW@���N8�?             5@        �       �                 pf�@      �?              @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �        	             *@        �       �                   @@@؇���X�?             @        �       �                   �@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 `�X#@�+Ĺ+�?6            �T@       �       �                   �:@�����?)            �O@       �       �                   �2@��?^�k�?            �A@        �       �                 ��Y @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     9@        �       �                   �;@�>4և��?             <@        ������������������������       �                      @        �       �                 �|�=@ȵHPS!�?             :@       �       �                 �|Y=@�X�<ݺ?             2@        ������������������������       �                     @        �       �                 ��) @�8��8��?	             (@       ������������������������       �                     $@        �       �                 �̜!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��)"@      �?              @       �       �                 @3�@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     *@        �       �                 �|�>@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��	0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     B@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������"iD��?&�-w���?iiiiii�?KKKKKK�?UUUUUU�?�������?              �?�$I�$I�?�m۶m��?              �?      �?        %I�$I��?n۶m۶�?      �?      �?              �?�������?�������?      �?      �?      �?                      �?              �?333333�?�������?UUUUUU�?�������?              �?�������?�������?              �?۶m۶m�?I�$I�$�?      �?      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?        �������?�������?      �?                      �?      �?                      �?�.�袋�?F]t�E�?      �?        �������?�������?              �?      �?        �c�!���?#8Q��4�?/�����?4և����?br1���?g���Q��?��+Q��?�]�ڕ��?�A�A�?|�W|�W�?              �?F]t�E�?]t�E]�?      �?                      �?]t�E�?/�袋.�?��y��y�?�0�0�?      �?      �?�B!��?���{��?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �������?�������?              �?      �?                      �?[��Z���?S+�R+��?�N��N��?�؉�؉�?1�0��?�y��y��?�;�;�?�؉�؉�?�$I�$I�?�m۶m��?              �?      �?        �������?UUUUUU�?              �?      �?        �{a���?a����?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?�؉�؉�?      �?                      �?333333�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?ى�؉��?�؉�؉�?      �?      �?      �?      �?      �?                      �?              �?      �?              �?        (ɟWY�?�ַC5�?t�E]t�?]t�E�?�{a���?��=���?Cy�5��?^Cy�5�?t�E]t�?]t�E�?      �?      �?�������?�������?              �?      �?      �?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?              �?      �?      �?      �?              �?      �?                      �?5H�4H��?�o��o��?�袋.��?]t�E�?333333�?�������?      �?        ۶m۶m�?�$I�$I�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        �?�������?;�;��?vb'vb'�?�������?�������?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?ى�؉��?�؉�؉�?F]t�E�?t�E]t�?      �?                      �?      �?              �?        �ذ��	�?�s�tD`�?      �?        �(ٵ���?%�6Q�k�?O���t:�?��b�X,�?�_FA@s�?���e�?      �?      �?]t�E�?t�E]t�?�������?333333�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?F]t�E�?t�E]t�?�q�q�?�q�q�?�������?�������?      �?              �?      �?              �?      �?              �?                      �?      �?        H�!��d�?x��m���?      �?        =
ףp=�?)\���(�?�D�a�Y�?���Id�?{�?g;�?4O��I�?      �?        ��.�?��6ͯ?              �?���c�?��N�©?���k(�?(�����?�%~F��?ہ�v`��?      �?        ��y��y�?�a�a�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        (፦ί�?���ˊ��?=��<���?�a�a�?_�_��?�A�A�?�������?�������?              �?      �?              �?        �$I�$I�?�m۶m��?              �?��N��N�?�؉�؉�?��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ6ޤhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������                           !@]@f�
�?�           8�@                                    @������?            �I@                                �-]@�X�<ݺ?             2@       ������������������������       �        	             .@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�q�q�?            �@@       	                           �?�GN�z�?             6@       
                           @$�q-�?             *@                                   @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@                                   @X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @                                   �?�eP*L��?             &@                                ��T?@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                    @և���X�?             @                               pf�@@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?               l                    �?�zv�X�?�           ��@               9                     @"pc�
�?�            @n@              $                     �?؀���˲?S            ``@                                  �H@ ����?)            @P@       ������������������������       �        "             L@                #                 ���I@�����H�?             "@        !       "                 ���;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        %       8                    �?�FVQ&�?*            �P@       &       '                 `f�)@�����?             E@        ������������������������       �                     &@        (       )                    �?��� ��?             ?@        ������������������������       �                     @        *       /                   �*@PN��T'�?             ;@        +       ,                    <@���Q��?             @        ������������������������       �                     �?        -       .                   �B@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        0       1                   �9@�C��2(�?             6@        ������������������������       �                     @        2       3                   �;@�r����?	             .@        ������������������������       �                     �?        4       5                   �E@@4և���?             ,@       ������������������������       �                     "@        6       7                    5@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     8@        :       O                    �?^H���+�?@            �[@        ;       @                   �-@�q��/��?            �H@        <       ?                    �?�q�q�?             @       =       >                   �+@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        A       N                 X�,A@���}<S�?             G@       B       K                    �?��S�ۿ?            �F@       C       D                 �|�6@��Y��]�?            �D@        ������������������������       �                     "@        E       J                    �?      �?             @@       F       G                 `fV&@XB���?             =@       ������������������������       �        	             1@        H       I                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        L       M                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        P       a                 ���1@�^�����?'             O@       Q       `                   @B@4�2%ޑ�?            �A@       R       _                    �?     ��?             @@       S       ^                    9@���B���?             :@       T       ]                   �7@      �?	             $@       U       Z                   �4@X�<ݚ�?             "@        V       Y                   �2@�q�q�?             @       W       X                 ��!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        [       \                 pff@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     @        ������������������������       �                     @        b       g                    @�>����?             ;@       c       f                 `fV6@ �q�q�?             8@        d       e                 ��)3@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        h       i                 ��T?@�q�q�?             @        ������������������������       �                     �?        j       k                   @D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        m       �                     �?��2(&�?            z@        n       }                 �|�<@x�(�3��?4            @S@        o       |                    �?X�Cc�?
             ,@       p       w                  �}S@�n_Y�K�?	             *@       q       r                    �?�<ݚ�?             "@        ������������������������       �                     @        s       t                   �;@�q�q�?             @        ������������������������       �                      @        u       v                 `f�D@      �?             @       ������������������������       �                      @        ������������������������       �                      @        x       y                 0�HU@      �?             @        ������������������������       �                      @        z       {                 ��)e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ~       �                 p�w@�<ݚ�?*            �O@              �                 `fF:@���*�?(             N@        ������������������������       �                     &@        �       �                    @@���c�H�?"            �H@        �       �                    �?     ��?             0@       �       �                 ���=@��S���?
             .@        �       �                    �?����X�?             @       �       �                 ���<@z�G�z�?             @        ������������������������       �                      @        �       �                 X��E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                  �>@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @       �       �                  �>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?<���D�?            �@@       �       �                  x;K@�J�4�?             9@        ������������������������       �                     .@        �       �                    �?���Q��?	             $@       �       �                 �U�T@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 03�M@      �?             @        ������������������������       �                     �?        �       �                 X��@@�q�q�?             @        ������������������������       �                     �?        �       �                    E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �C@�hQ����?�            Pu@       �       �                 ��@(71����?�            �r@        �       �                    �?hA� �?,            �Q@        �       �                 ���@R���Q�?             4@        �       �                 �|�9@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �5@z�G�z�?             $@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|=@      �?              @        ������������������������       �                     @        �       �                 �|�=@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     I@        �       �                 ��`3@����/�?�            `l@       �       �                 ��d2@�MI8d�?r             g@       �       �                   @C@R���Q�?p            �f@       �       �                    �?T���D9�?n            �e@        �       �                    �?ҳ�wY;�?             1@       �       �                 �|Y=@������?
             .@        �       �                   �1@�q�q�?             @        ������������������������       �                      @        �       �                     @      �?             @        ������������������������       �                     �?        �       �                 ��Y&@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        �       �                 �|�=@���1���?b            �c@       �       �                    �?P���Q�?K             ^@        ������������������������       �                     @        �       �                    �?P���Q�?G            �\@       �       �                     @�}�+r��?F            �\@        ������������������������       �                     &@        �       �                 �?$@p�eU}�??            �Y@        ������������������������       �      �?             @        �       �                   �0@Pa�	�?=            �X@        �       �                 pFD!@؇���X�?             @        ������������������������       �      �?             @        ������������������������       �                     @        �       �                 �?�@��<b�ƥ?8             W@        ������������������������       �                    �G@        �       �                 @3�@`Ӹ����?             �F@        �       �                   �4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 pf� @��Y��]�?            �D@        �       �                 ��) @P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     �?        �       �                     @p9W��S�?             C@        �       �                 `fF)@r�q��?             (@        ������������������������       �                     @        �       �                    @@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �&B@$��m��?             :@        ������������������������       �                     @        �       �                 @3�@8�A�0��?             6@        �       �                    A@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                 ���!@d}h���?             ,@        ������������������������       �                     @        �       �                 ��)@և���X�?             @        �       �                   �?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     @z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �2@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �?@�Ń��̧?             E@       ������������������������       �                     =@        �       �                     @$�q-�?	             *@        ������������������������       �                     @        �       �                 �T�E@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     F@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������ߺ?9���?C����v�?�?xxxxxx�?�q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?]t�E�?�袋.��?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?r�q��?      �?                      �?t�E]t�?]t�E�?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?                      �?��.���?�袋.��?F]t�E�?/�袋.�?�i��?h�T��? �����? �����?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?|���?>����?�a�a�?=��<���?              �?�B!��?�{����?              �?h/�����?&���^B�?�������?333333�?      �?              �?      �?              �?      �?        F]t�E�?]t�E�?              �?�?�������?      �?        �$I�$I�?n۶m۶�?              �?�������?�������?              �?      �?                      �?�g�`�|�?L�Ϻ��?և���X�?/����?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        d!Y�B�?ӛ���7�?�?�������?������?8��18�?              �?      �?      �?�{a���?GX�i���?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?              �?        !�B�?���{��?�A�A�?�������?      �?      �?ى�؉��?��؉���?      �?      �?�q�q�?r�q��?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?      �?              �?      �?              �?                      �?              �?      �?        �Kh/��?h/�����?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ��.���?t�E]t�?(�Y�	q�?�wL��?�m۶m��?%I�$I��?ى�؉��?;�;��?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?                      �?9��8���?�q�q�?""""""�?wwwwww�?      �?        4և����?/�����?      �?      �?�?�������?�m۶m��?�$I�$I�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?              �?      �?              �?333333�?�������?      �?      �?      �?                      �?      �?              �?        |���?|���?�z�G��?{�G�z�?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?�<��3��?�f�a��?�F�1V�?��pN�?���?_�_�?333333�?333333�?�������?�������?              �?      �?        �������?�������?      �?      �?              �?      �?              �?      �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?        L���D��?҂��z�?��L���?L�Ϻ��?333333�?333333�?���NV��?��Ħ��?�������?�������?wwwwww�?�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�3���?7a~W��?ffffff�?�������?      �?        �ø_�T�?��s���?�5��P�?(�����?      �?        (�J��"�?��VCӭ?      �?      �?|���?|���?۶m۶m�?�$I�$I�?      �?      �?      �?        ��7��M�?d!Y�B�?      �?        ?�>��?l�l��?      �?      �?              �?      �?        8��18�?������?ffffff�?�������?      �?                      �?      �?              �?        �k(����?l(�����?�������?UUUUUU�?      �?        333333�?�������?      �?                      �?�N��N��?vb'vb'�?      �?        颋.���?/�袋.�?      �?      �?              �?      �?        I�$I�$�?۶m۶m�?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?              �?        �������?�������?      �?                      �?�������?333333�?      �?                      �?��<��<�?�a�a�?      �?        �؉�؉�?;�;��?      �?              �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��{hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       ^                    �?ʡ�;S��?�           8�@               #                    �?0,Tg��?�            �o@                                  �-@L������?1            @R@                                P��+@�q�q�?             @        ������������������������       �                     @                                   @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        	                        ��.@�qM�R��?,            �P@        
                           �?��<b���?             7@                                  �7@���Q��?             @        ������������������������       �                     �?                                �|Y=@      �?             @        ������������������������       �                     �?                                ��%@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                    @�����H�?             2@        ������������������������       �                     @                                   �?�r����?
             .@                               �|�9@@4և���?	             ,@        ������������������������       �                     @                                 ��@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?               "                    �?`���i��?             F@              !                     �?      �?             @@                                 �H@`2U0*��?             9@       ������������������������       �                     6@                                 83F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        $       M                 �|�=@��bu<	�?j            `f@       %       F                    �?�5g����?A            @[@       &       '                     @�lg����?2            �U@        ������������������������       �                    �@@        (       +                 pf�@Fmq��?            �J@        )       *                 �|Y:@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ,       A                    �?v�X��?             F@       -       6                 @3�@������?             >@        .       1                 �&B@�eP*L��?             &@        /       0                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        2       3                 P�@���Q��?             @        ������������������������       �                      @        4       5                   �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        7       8                  �#@�S����?             3@        ������������������������       �                      @        9       :                    '@���!pc�?             &@        ������������������������       �                     �?        ;       @                 �|�;@z�G�z�?             $@       <       ?                    4@�����H�?             "@       =       >                 `F�+@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        B       E                   �;@X�Cc�?	             ,@       C       D                 @3�2@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        G       H                     @
;&����?             7@        ������������������������       �                     @        I       L                 �|�:@      �?
             0@       J       K                    *@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        N       Y                     @z�G�z�?)            �Q@       O       R                   �'@,�+�C�?!            �K@        P       Q                   �J@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        S       T                   �E@@9G��?            �H@       ������������������������       �                     @@        U       X                    :@�t����?             1@        V       W                  ��9@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        Z       ]                    �?�q�q�?             .@        [       \                   �>@      �?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        _       �                     �?"~��F��?           �|@        `       �                    K@�&!��?8            �U@       a       z                   �B@� �	��?/            �R@        b       y                   @G@^������?            �A@       c       d                 ��I/@�q�����?             9@        ������������������������       �                     @        e       x                   @>@�����?             3@       f       g                 03k:@և���X�?             ,@        ������������������������       �                      @        h       o                    �?      �?
             (@        i       n                    �?�q�q�?             @       j       m                 �ܵ<@z�G�z�?             @        k       l                 ��";@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        p       q                   �<@�q�q�?             @        ������������������������       �                     �?        r       s                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        t       w                 X��B@      �?             @       u       v                 `fF<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        {       �                    H@      �?             D@       |       }                    &@     ��?             @@        ������������������������       �                     �?        ~       �                    �?��� ��?             ?@              �                 03�S@$�q-�?             :@       ������������������������       �        
             ,@        �       �                 X��@@r�q��?             (@       ������������������������       �                      @        �       �                   �D@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    9@���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @       �       �                   �?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �H@      �?              @        ������������������������       �                     @        �       �                   @I@      �?             @       �       �                 `f^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�C��2(�?	             &@        ������������������������       �                     @        �       �                   �R@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @X/I2w��?�            Pw@        �       �                    @b�2�tk�?             2@       �       �                   �C@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��	}g�?�            0v@        �       �                 ��K.@R���Q�?             D@       �       �                     @�r����?             >@        ������������������������       �                     @        �       �                 pF�#@�J�4�?             9@       �       �                 �� @�LQ�1	�?             7@       �       �                   �6@؇���X�?             5@        ������������������������       �                     �?        �       �                 ���@ףp=
�?             4@        ������������������������       �                     @        �       �                   @@8�Z$���?             *@        �       �                 �|=@      �?              @        ������������������������       �                     @        ������������������������       �      �?              @        �       �                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    /@      �?             $@        ������������������������       �                      @        �       �                 м;4@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                     @,B�r��?�            �s@        �       �                   �@@Pa�	�?%            �P@       ������������������������       �                     A@        �       �                   �*@      �?             @@        �       �                 `f�)@8�Z$���?             *@        ������������������������       �                     @        �       �                   �A@����X�?             @        ������������������������       �                     �?        �       �                   �C@r�q��?             @        ������������������������       �                     @        �       �                    G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        �       �                   �>@�cX1!��?�             o@       �       �                    �?�7��?t            `h@        ������������������������       �                    �A@        �       �                    $@      �?_             d@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                 `f�9@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �T�I@��}� �?[            `c@       �       �                   �:@���	���?X            �b@       �       �                    �?(;L]n�?5            �V@       �       �                   �4@@�)�n�?0            @U@       �       �                   �1@��p\�?            �D@        ������������������������       �                     (@        �       �                   �2@ܷ��?��?             =@        �       �                 ��Y @      �?             @       �       �                  s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 0S5 @HP�s��?             9@       �       �                 �?�@r�q��?             (@       ������������������������       �                      @        �       �                   �3@      �?             @        ������������������������       �      �?              @        ������������������������       �      �?              @        ������������������������       �                     *@        ������������������������       �                     F@        ������������������������       �                     @        �       �                 ��) @��GEI_�?#            �N@       ������������������������       �                     I@        �       �                   �;@���|���?	             &@        ������������������������       �                      @        �       �                 pf� @�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                 p�O@      �?             @       �       �                    ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �                          �?�+$�jP�?             K@       �       �                    �?��[�p�?            �G@        ������������������������       �                     �?        �                       �T)D@��<b���?             G@       �       �                 �&B@,���i�?            �D@        ������������������������       �                     4@        �       �                   �?@���N8�?             5@        ������������������������       �                     �?        �                        @3�@z�G�z�?             4@        �       �                 �?�@X�<ݚ�?             "@       �       �                    A@r�q��?             @        �       �                   �@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������N���I5�?d�~`l��?1�0��?�y��y��?����?�Ǐ?~�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?        ���@��?�n�Wc"�?��Moz��?��,d!�?333333�?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?              �?�?�������?�$I�$I�?n۶m۶�?              �?�������?�������?      �?                      �?      �?        F]t�E�?F]t�E�?      �?      �?{�G�z�?���Q��?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?��49ȼ�?��e㛡�?\������?R1�:#�?�}A_��?}A_��?              �?�x+�R�?~�	�[�?�q�q�?�q�q�?              �?      �?        �.�袋�?颋.���?wwwwww�?�?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?(������?^Cy�5�?      �?        F]t�E�?t�E]t�?              �?�������?�������?�q�q�?�q�q�?�������?�������?              �?      �?              �?                      �?%I�$I��?�m۶m��?UUUUUU�?�������?              �?      �?              �?        Y�B��?�Mozӛ�?              �?      �?      �?r�q��?�q�q�?      �?                      �?      �?        �������?�������?��)A��?�}��7��?UUUUUU�?UUUUUU�?              �?      �?        9/���?������?              �?�?<<<<<<�?�������?333333�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        �A^%���?���j�1�?֔5eMY�?S֔5eM�?�Q����?)\���(�?_�_��?uPuP�?���Q��?�p=
ף�?      �?        ^Cy�5�?Q^Cy��?۶m۶m�?�$I�$I�?              �?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?      �?      �?      �?      �?              �?�{����?�B!��?�؉�؉�?;�;��?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?        333333�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?u>q��e�?[v�cӼ?9��8���?�8��8��?]t�E]�?F]t�E�?              �?      �?                      �?��j�4�?(�/��Z�?�������?�������?�������?�?      �?        �z�G��?{�G�z�?��Moz��?Y�B��?۶m۶m�?�$I�$I�?              �?�������?�������?      �?        ;�;��?;�;��?      �?      �?      �?              �?      �?�������?�������?              �?      �?              �?              �?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?        >��=���?��?|���?|���?      �?              �?      �?;�;��?;�;��?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?        I�dn�?��ٌ?��[��[�?�A�A�?      �?              �?      �?�������?�������?      �?              �?      �?              �?      �?        $^E�U$�?��ۡ��?�z=��?��^x/��?�������?�?�������?�?�]�ڕ��?��+Q��?      �?        ��=���?a���{�?      �?      �?      �?      �?      �?                      �?      �?        q=
ףp�?{�G�z�?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?      �?      �?              �?              �?        �d����?;ڼOqɰ?      �?        ]t�E]�?F]t�E�?              �?9��8���?�q�q�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        /�����?B{	�%��?�
br1�?m�w6�;�?      �?        ��,d!�?��Moz��?�����?8��18�?      �?        �a�a�?��y��y�?              �?�������?�������?r�q��?�q�q�?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ?{�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM	hjh))��}�(h,h/h0M	��h2h3h4hph<�h=Kub������       v                     @>AU`�z�?�           8�@               !                    �?�p����?�            Pt@                                  �8@���j��?7             W@                                   �?PN��T'�?             ;@       ������������������������       �                     3@                                ���Q@      �?              @        ������������������������       �                     @        ������������������������       �                     @        	       
                    �?�4��?&            @P@        ������������������������       �                     ?@                                 p�w@ҳ�wY;�?             A@                               �ܵ<@>���Rp�?             =@        ������������������������       �                     @                                 	>@ �o_��?             9@                                ���=@      �?             @                               X��E@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                 �>@��s����?             5@        ������������������������       �                      @                                p"�X@�	j*D�?
             *@                                   �?X�<ݚ�?             "@                               x�R@      �?              @                               X�lA@�q�q�?             @        ������������������������       �                     @                                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        "       i                    �?�=�Ȇ��?�             m@       #       J                     �?�-��ē�?o            �e@        $       %                    �?�\��N��?1             S@        ������������������������       �                     8@        &       9                  i?@�	j*D�?!             J@        '       (                   �<@
j*D>�?             :@        ������������������������       �                     @        )       8                   @>@�LQ�1	�?             7@       *       +                 ��$:@����X�?             5@        ������������������������       �                     @        ,       7                    R@ҳ�wY;�?	             1@       -       0                    D@������?             .@        .       /                 `fF<@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        1       6                 `f�;@ףp=
�?             $@       2       3                   @G@؇���X�?             @        ������������������������       �                     @        4       5                    J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        :       =                  x#J@���B���?             :@        ;       <                 �|�<@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        >       ?                 `�iJ@�q�q�?
             (@        ������������������������       �                      @        @       G                 03�U@z�G�z�?	             $@       A       F                   @K@      �?              @        B       C                    7@      �?             @        ������������������������       �                      @        D       E                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        H       I                 �w|c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        K       d                   �E@uvI��?>            �X@       L       Y                    �?�L"p�?3            �T@        M       X                   �7@�8��8��?             B@       N       O                   �;@@�0�!��?             1@        ������������������������       �                      @        P       Q                 `f�)@��S�ۿ?             .@        ������������������������       �                     @        R       W                   �,@�����H�?             "@       S       T                   �B@؇���X�?             @       ������������������������       �                     @        U       V                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     3@        Z       c                    1@=QcG��?            �G@       [       b                   �C@     ��?             @@       \       a                    &@h�����?             <@        ]       ^                    @@4և���?	             ,@        ������������������������       �                     @        _       `                    5@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        
             ,@        ������������������������       �      �?             @        ������������������������       �        	             .@        e       h                 `f'@��S�ۿ?             .@        f       g                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             &@        j       u                   �L@�:�B��?(            �M@       k       r                    <@�NW���?%            �J@       l       q                    �?�?�|�?            �B@       m       p                    @(;L]n�?             >@        n       o                 ��1V@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     9@        ������������������������       �                     @        s       t                    �?     ��?             0@       ������������������������       �        
             *@        ������������������������       �                     @        ������������������������       �                     @        w                         �C@vp�*�?�             x@       x                          @zoB����?�            �u@       y       �                    �?`��b�?�            �u@        z       �                 ���@z�H}��?C            �Z@        {       ~                    �?��� ��?             ?@        |       }                 0��@      �?             @       ������������������������       �                     @        ������������������������       �                     @               �                    �?`2U0*��?             9@       �       �                 ���@���7�?             6@       �       �                 03S@�C��2(�?             &@        ������������������������       �                     @        �       �                 �|�9@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        �       �                   0:@      �?1             S@       �       �                 �|Y=@)O���?/             R@        �       �                 �&�)@�t����?             1@        ������������������������       �                      @        �       �                    �?X�<ݚ�?             "@       �       �                    �?      �?              @       �       �                 �0@���Q��?             @       �       �                    �?      �?             @       �       �                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?\�����?!            �K@        �       �                    �?�q�q�?             8@       ������������������������       �                     3@        ������������������������       �                     @        �       �                 �?$'@��a�n`�?             ?@       �       �                 ��(@      �?             8@       �       �                  s�@�S����?	             3@        ������������������������       �                     �?        ������������������������       �r�q��?             2@        ������������������������       �                     @        �       �                    �?և���X�?             @       �       �                  �v6@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�B+w@�?�            �m@        �       �                   @1@�ՙ/�?&            �O@       �       �                    �?Hث3���?            �C@       �       �                 ���@)O���?             B@        �       �                  s@�<ݚ�?             "@        ������������������������       �                      @        �       �                 pff@����X�?             @       �       �                 �|Y:@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �|�=@��}*_��?             ;@       �       �                   �3@�GN�z�?             6@        �       �                    �?z�G�z�?             @       �       �                 �&B@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �@�IєX�?
             1@        �       �                 �&B@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��p@@r�q��?             8@       �       �                    �?�<ݚ�?             2@        ������������������������       �                     @        �       �                    @�	j*D�?
             *@        ������������������������       �                      @        �       �                   �>@"pc�
�?	             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        �       �                    )@x̓��s�?t            �e@        �       �                 `f�7@      �?             $@        ������������������������       �                     @        ������������������������       �                     @        �                         @C@,�+�C�?m            �d@       �                          �?��M6�?k            `d@       �       �                 �?�@�E����?g            �c@        �       �                   �7@�?�|�?2            �R@        ������������������������       �                     A@        �       �                   �8@P���Q�?             D@        �       �                   �@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|Y=@�?�|�?            �B@        ������������������������       �                     1@        �       �                  sW@P���Q�?             4@        �       �                 �|Y?@؇���X�?             @       �       �                 pf�@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �        
             *@        �       �                   �2@��Lɿ��?5            �T@        �       �                   �1@      �?              @       ������������������������       �                     @        �       �                 ��Y @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 @3�@���Lͩ�?0            �R@        �       �                   �=@�q�q�?             @        ������������������������       �                      @        �       �                   �?@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 ��) @D��*�4�?+            @Q@        ������������������������       �                     5@        �       �                 ��y @8��8���?             H@        ������������������������       �                     �?        �                        �|Y=@dP-���?            �G@       �       �                 �T)D@��� ��?             ?@       �       �                    (@ �Cc}�?             <@       �       �                 ���"@@�0�!��?	             1@       �       �                   �:@�����H�?             "@       ������������������������       �                     @        �       �                    <@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �<@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        �       �                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     @                              ��	0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                @C@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �B@        �*       h�h))��}�(h,h/h0M	KK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?�<�@�0�?�a�ߔ��?!Y�B�?ozӛ���?h/�����?&���^B�?              �?      �?      �?              �?      �?        �Z��Z��?�R+�R+�?              �?�������?�������?�i��F�?GX�i���?      �?        
ףp=
�?�Q����?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?z��y���?�a�a�?      �?        vb'vb'�?;�;��?r�q��?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?                      �?���c�?p�2N�?�l����?A&�dR�?�5��P�?y�5���?              �?vb'vb'�?;�;��?b'vb'v�?;�;��?              �?Nozӛ��?d!Y�B�?�m۶m��?�$I�$I�?      �?        �������?�������?wwwwww�?�?�������?333333�?              �?      �?        �������?�������?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?                      �?              �?��؉���?ى�؉��?n۶m۶�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?      �?      �?      �?              �?      �?              �?      �?              �?              �?      �?              �?      �?        ��X��?
^N��)�?�FS���?rY1P��?UUUUUU�?UUUUUU�?�������?ZZZZZZ�?      �?        �?�������?              �?�q�q�?�q�q�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?x6�;��?AL� &W�?      �?      �?�m۶m��?�$I�$I�?n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?              �?              �?      �?      �?        �������?�?      �?      �?              �?      �?              �?        �pR���?�c+����?�x+�R�?萚`���?к����?*�Y7�"�?�?�������?�������?�������?              �?      �?                      �?              �?      �?      �?              �?      �?              �?        �~����?c�z���?xJW�?"��ע��?���+M�?��P��?�S�rp�?��XQ�?�{����?�B!��?      �?      �?              �?      �?        ���Q��?{�G�z�?�.�袋�?F]t�E�?]t�E�?F]t�E�?      �?        �������?UUUUUU�?              �?      �?              �?              �?              �?      �?��8��8�?9��8���?�������?�������?              �?r�q��?�q�q�?      �?      �?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?߰�k��?A��)A�?�������?UUUUUU�?              �?      �?        �c�1��?�s�9��?      �?      �?(������?^Cy�5�?      �?        �������?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?      �?        ��|��|�?V�V��?�<��<��?�a�a�?��-��-�?�i�i�?9��8���?��8��8�?�q�q�?9��8���?              �?�$I�$I�?�m۶m��?�������?333333�?              �?      �?                      �?_B{	�%�?B{	�%��?�袋.��?]t�E�?�������?�������?      �?      �?      �?                      �?              �?�?�?      �?      �?      �?                      �?      �?                      �?              �?�������?UUUUUU�?9��8���?�q�q�?      �?        vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?      �?                      �?      �?        v��4��?L�w�Z޸?      �?      �?              �?      �?        �}��7��?��)A��?��g*��?|��¬F�?�}��	��?�����?*�Y7�"�?к����?      �?        ffffff�?�������?UUUUUU�?UUUUUU�?              �?      �?        *�Y7�"�?к����?      �?        ffffff�?�������?۶m۶m�?�$I�$I�?�������?�������?      �?              �?      �?      �?              �?        �������?rY1P»?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �6�i�?�K~��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ہ�v`��?)�3J���?      �?        �������?�������?              �?�����F�?W�+�ɵ?�{����?�B!��?%I�$I��?۶m۶m�?ZZZZZZ�?�������?�q�q�?�q�q�?      �?        �������?�������?              �?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?      �?              �?      �?              �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��}whG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       V                    �?"��p�?�           8�@               G                   �?@&j���$�?�             o@              2                    �?�{����?k             f@              1                 м�9@�('+��?T            �a@                                 �,@�Sb(�	�?=             [@        ������������������������       �                     (@                                �B,@r�q��?5             X@              	                    �?<ݚ�?(             R@        ������������������������       �                     =@        
                            @�&!��?            �E@        ������������������������       �                     (@                                  �3@`՟�G��?             ?@                                �&B@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                pff@��H�}�?             9@                                pff@����X�?             @                                ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �7@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  �&@�<ݚ�?             2@                               @3�@      �?	             0@                                  �9@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @                                   �-@      �?             8@        ������������������������       �                     @        !       (                 ��1@�����?             3@        "       %                    �?X�<ݚ�?             "@        #       $                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        &       '                 �|�<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        )       *                   �;@z�G�z�?             $@        ������������������������       �                     @        +       ,                 �|�<@�q�q�?             @        ������������������������       �                     �?        -       .                 �|Y>@z�G�z�?             @        ������������������������       �                      @        /       0                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �A@        3       8                    �?j���� �?             A@        4       7                 ��Ya@z�G�z�?             @        5       6                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        9       F                    @П[;U��?             =@       :       ?                     @���>4��?             <@       ;       <                 ��[@d}h���?
             ,@       ������������������������       �                     @        =       >                 Ъ�c@      �?              @        ������������������������       �                     @        ������������������������       �                     @        @       A                    @����X�?             ,@        ������������������������       �                      @        B       E                 �|�:@r�q��?             (@       C       D                 ��L6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        H       Q                     @4?,R��?-             R@       I       J                     �?P����?%            �M@       ������������������������       �                    �B@        K       L                   �B@���7�?             6@       ������������������������       �                     *@        M       P                    �?�����H�?             "@       N       O                    D@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        R       U                   �5@�	j*D�?             *@        S       T                   �A@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        W                           �?I����?           �|@       X       �                    �?Ry���?           �z@        Y       n                 �|Y=@�!���?.             Q@        Z       a                 �&�)@r�q��?             8@        [       `                   @@      �?             (@       \       _                    �?և���X�?             @       ]       ^                   �7@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        b       c                    3@�q�q�?
             (@        ������������������������       �                     @        d       m                    �?      �?              @       e       f                 ���0@և���X�?             @        ������������������������       �                      @        g       l                     @���Q��?             @       h       k                     �?      �?             @       i       j                   �8@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        o       �                 p�w@�������?             F@       p       }                     �?r�q��?             E@        q       |                 �UkT@���y4F�?             3@       r       {                   �J@�q�q�?             (@       s       t                 ���<@      �?              @        ������������������������       �                     �?        u       z                    �?և���X�?             @       v       y                 X��C@�q�q�?             @       w       x                 ��2>@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ~       �                    �?�LQ�1	�?             7@              �                   @@�C��2(�?             6@       �       �                 ���@r�q��?             (@        ������������������������       �                     @        �       �                 �|�=@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @�2��g�?�            �v@        �       �                    �?���Q��?             $@        ������������������������       �                      @        �       �                   l@@      �?              @       �       �                 ��|2@؇���X�?             @        ������������������������       �                     @        �       �                 ���7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                     �?\��0���?�            v@        �       �                  x#J@
��[��?&            @P@       �       �                   �<@���c�H�?            �H@        �       �                   �;@����X�?             @        ������������������������       �                     �?        �       �                 `f�D@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    R@؇���X�?             E@       �       �                   �>@ףp=
�?             D@       �       �                   @>@���y4F�?             3@       �       �                 03k:@�t����?             1@        �       �                   �9@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �C@@4և���?             ,@        �       �                 �|�?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �        
             5@        ������������������������       �                      @        �       �                 �|Y<@     ��?             0@        �       �                    7@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���!pc�?	             &@       �       �                    �?և���X�?             @        ������������������������       �                     �?        �       �                 `�iJ@      �?             @        ������������������������       �                     �?        �       �                   �B@���Q��?             @        ������������������������       �                      @        �       �                 ��<R@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �2@�5?,R�?�             r@        �       �                 ��Y @"pc�
�?            �@@        �       �                 ��@�q�q�?             "@        ������������������������       �                      @        �       �                    1@؇���X�?             @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     8@        �       �                 0��G@�:�]��?�            �o@       �       �                 ���@0{�v��?�            @o@        ������������������������       �                    �H@        �       �                   �<@�qM�R��?}             i@        �       �                 @3�!@��ɉ�?+            @P@       �       �                   � @ �#�Ѵ�?            �E@       �       �                   �4@ ���J��?            �C@        �       �                 @3�@�C��2(�?             &@       �       �                 �?�@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     <@        �       �                   �:@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     6@        �       �                     @�t����?R             a@        �       �                 `f�)@�nkK�?             G@        ������������������������       �        	             0@        �       �                    �?��S�ۿ?             >@       �       �                    C@HP�s��?             9@        ������������������������       �                     &@        �       �                    ,@؇���X�?             ,@        �       �                   �F@      �?              @        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|Y=@���V��?9            �V@        �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                   `!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?���H��?6             U@       �       �                    �?,���i�?4            �T@        �       �                 ��(@ ��WV�?             :@       �       �                 X�I@P���Q�?
             4@       ������������������������       ��}�+r��?	             3@        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �?@�X�C�?'             L@       �       �                 �|�=@�'�`d�?            �@@       �       �                  sW@؇���X�?             <@        ������������������������       ����Q��?             @        �       �                 ��) @�nkK�?             7@       ������������������������       �                     0@        �       �                 pf� @؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 @3�@���}<S�?             7@        �       �                   @C@      �?              @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �        
             .@        ������������������������       �                      @        �       �                    ;@���Q��?             @        ������������������������       �                     �?        �       �                 �|�>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                 �?�g�y��?             ?@                                  �?      �?              @                               "&d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 *@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        	                         @�û��|�?             7@       
                          �?8�A�0��?             6@        ������������������������       �                      @                                 #@��Q��?             4@                              pf�C@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������J54v��?l�����?ְ�"NT�?��Bw�j�?�Br���?��F($�?����#T�?R��*�?�Kh/���?�Kh/��?              �?UUUUUU�?UUUUUU�?��8��8�?�q�q�?              �?S֔5eM�?֔5eMY�?              �?�1�c��?�s�9��?UUUUUU�?�������?      �?                      �?{�G�z�?
ףp=
�?�$I�$I�?�m۶m��?      �?      �?              �?      �?        �������?�������?              �?      �?        9��8���?�q�q�?      �?      �?�m۶m��?�$I�$I�?      �?                      �?      �?                      �?      �?      �?      �?        Q^Cy��?^Cy�5�?r�q��?�q�q�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?ZZZZZZ�?�������?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?��=���?�{a���?n۶m۶�?I�$I�$�?۶m۶m�?I�$I�$�?              �?      �?      �?      �?                      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?r�q��?�8��8��?'u_[�?�V'u�?              �?F]t�E�?�.�袋�?              �?�q�q�?�q�q�?�$I�$I�?۶m۶m�?      �?                      �?              �?vb'vb'�?;�;��?      �?      �?              �?      �?              �?        g�'�Y��?dj`��?U�����?��0b�?�������?�������?UUUUUU�?UUUUUU�?      �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?�$I�$I�?۶m۶m�?      �?        �������?333333�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?t�E]t�?/�袋.�?�������?UUUUUU�?6��P^C�?(������?UUUUUU�?UUUUUU�?      �?      �?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?�������?333333�?              �?      �?                      �?      �?              �?              �?        ��Moz��?Y�B��?]t�E�?F]t�E�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?              �?                      �?              �?;G����?㺥��?�������?333333�?      �?              �?      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        @����?�:��?7r#7r#�?�����?4և����?/�����?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?�$I�$I�?�������?�������?6��P^C�?(������?<<<<<<�?�?UUUUUU�?UUUUUU�?      �?                      �?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?                      �?      �?      �?�������?�������?      �?                      �?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?              �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?�q�q�?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?        }}}}}}�?�?V-��?;�O��n�?      �?        �n�Wc"�?���@��??�?��? �����?�/����?�}A_Ч?��-��-�?�A�A�?]t�E�?F]t�E�?�������?�������?      �?              �?      �?      �?              �?              �?      �?      �?                      �?      �?        <<<<<<�?�?�Mozӛ�?d!Y�B�?      �?        �������?�?q=
ףp�?{�G�z�?      �?        ۶m۶m�?�$I�$I�?      �?      �?333333�?�������?      �?              �?              �?        [�[��?�>�>��?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�0�0�?��y��y�?�����?8��18�?O��N���?;�;��?ffffff�?�������?�5��P�?(�����?      �?              �?        �m۶m��?%I�$I��?6�d�M6�?'�l��&�?۶m۶m�?�$I�$I�?�������?333333�?�Mozӛ�?d!Y�B�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        �������?333333�?      �?                      �?ӛ���7�?d!Y�B�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?        333333�?�������?              �?      �?      �?      �?                      �?�B!��?��{���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?        8��Moz�?��,d!�?颋.���?/�袋.�?              �?�������?ffffff�?�q�q�?9��8���?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�,�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM)hjh))��}�(h,h/h0M)��h2h3h4hph<�h=Kub������                       `f~I@���$ӡ�?�           8�@              [                     @��n:���?x           ��@               &                 �J+@�5�uԞ�?z            @i@               	                    �?������?.             Q@                                ��Y(@�q�q�?             @        ������������������������       �                     �?                                X��E@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        
       %                    �?�n`���?+             O@                                  �?`��:�?*            �N@                                  �:@���Q��?             .@        ������������������������       �                      @                                  �J@�	j*D�?
             *@                                 �B@"pc�
�?	             &@        ������������������������       �                     @                                   D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                   4@���.�6�?             G@                                  �2@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                `fF)@���N8�?             E@       ������������������������       �                     5@               $                   �*@�����?             5@                                  @@�t����?
             1@        ������������������������       �                     @                                  �A@r�q��?             (@        ������������������������       �      �?              @                #                    G@ףp=
�?             $@       !       "                   �C@r�q��?             @        ������������������������       �                     �?        ������������������������       �z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        '       0                    �?��:c���?L            �`@        (       )                  ��9@����?�?            �F@        ������������������������       �        
             3@        *       /                    :@ ��WV�?             :@        +       .                    �?ףp=
�?             $@       ,       -                    D@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             0@        1       6                 `ff:@:��?2            @V@        2       3                     �?�r����?             >@        ������������������������       �                      @        4       5                    "@؇���X�?             <@        ������������������������       �                     @        ������������������������       �                     8@        7       Z                 �D B@TV����?!            �M@       8       9                   �<@Rg��J��?            �H@        ������������������������       �                     $@        :       E                    �?�e����?            �C@        ;       @                   @@@�q�q�?             (@        <       ?                 �|�=@z�G�z�?             @       =       >                 ��2>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        A       B                    <@؇���X�?             @        ������������������������       �                     @        C       D                   �H@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        F       Y                   �Q@�q�q�?             ;@       G       X                  i?@�	j*D�?             :@       H       W                   @>@�ՙ/�?             5@       I       V                     �?�E��ӭ�?             2@       J       K                 �|Y=@     ��?	             0@        ������������������������       �                     @        L       U                   �J@�n_Y�K�?             *@       M       T                 `fF<@      �?             $@       N       S                    H@      �?              @       O       P                 �|�?@����X�?             @        ������������������������       �                      @        Q       R                   �C@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        \       �                    �?H��%�R�?�            �x@        ]       �                 ��Y7@�qs�_�?M            �Z@       ^       e                 ��@��p �?;            �T@        _       `                  �[@���}<S�?             7@        ������������������������       �                     @        a       d                    �?�t����?             1@       b       c                 P�@      �?             0@        ������������������������       �                     �?        ������������������������       �        
             .@        ������������������������       �                     �?        f       g                    @Ɣ��Hr�?+            �M@        ������������������������       �                     @        h       �                  �2@���3L�?'             K@       i       �                 ���1@z�J��?#            �G@       j       y                   �9@v�2t5�?             �D@        k       v                    �?b�2�tk�?             2@       l       q                   �3@���Q��?             .@        m       n                    �?r�q��?             @        ������������������������       �                     @        o       p                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        r       u                 pff@�����H�?             "@        s       t                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        w       x                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        z       �                    �?��+7��?             7@       {       |                 @3�@      �?             4@        ������������������������       �                     @        }       ~                    �?�t����?             1@        ������������������������       �                     �?               �                   �:@      �?             0@        ������������������������       �                     �?        �       �                    �?z�G�z�?             .@       �       �                   �D@"pc�
�?	             &@       �       �                 �|Y>@ףp=
�?             $@       �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                 pf&(@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �&@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @�J�4�?             9@       �       �                  ��8@P���Q�?             4@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        �       �                 ��A>@���Q��?             @        ������������������������       �                     �?        �       �                   @D@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?\�ih�<�?�            �q@        �       �                 03�-@�G�z�?             D@       �       �                 �&�)@r٣����?            �@@       �       �                 �y�#@������?             >@       �       �                 �-!@d}h���?             <@       �       �                   �6@�+e�X�?             9@        �       �                   �2@z�G�z�?             @        �       �                 ��}@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���@ףp=
�?             4@        ������������������������       �                      @        �       �                 �|�=@r�q��?             (@       �       �                   @@�<ݚ�?             "@       �       �                 �|�:@      �?              @        ������������������������       �                     �?        ������������������������       �����X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    /@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    #@`U���H�?�            �n@        �       �                    �?��.k���?	             1@       �       �                    �?�q�q�?             "@        ������������������������       �                     @        �       �                 03�;@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 pf�C@      �?              @       �       �                    @r�q��?             @       �       �                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���@�˹�m��?�            �l@        ������������������������       �                     8@        �       �                    �?l��\��?            �i@        �       �                   `3@�t����?             A@       �       �                  ��@��a�n`�?             ?@        ������������������������       �                      @        �       �                 ��(@�LQ�1	�?             7@       �       �                 �|Y=@     ��?             0@        ������������������������       �                     �?        �       �                 X�I@�r����?
             .@       ������������������������       �8�Z$���?	             *@        ������������������������       �                      @        ������������������������       �                     @        �       �                 03�7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ���@�m(�X�?k            @e@        ������������������������       �                     @        �                       `f�'@��
�π�?j            �d@       �       �                 �|�=@���D�k�?S            �`@       �       �                   �0@p�qG�?<             X@        �       �                 pf�@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        �       �                 �?�@�nkK�?9             W@       �       �                 �|�<@@��8��?             H@       ������������������������       �                     >@        �       �                  sW@�X�<ݺ?             2@        �       �                 ��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     .@        �       �                 @3�@t��ճC�?             F@        �       �                   �4@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 ��) @�7��?            �C@        ������������������������       �                     *@        �       �                 0SE @$�q-�?             :@        ������������������������       �                     �?        �       �                 @3�!@`2U0*��?             9@       �       �                 pf� @��S�ۿ?	             .@        ������������������������       �                     @        �       �                   �:@�8��8��?             (@       ������������������������       �                     $@        �       �                 �|Y<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �?@�MI8d�?            �B@        �       �                 �?�@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �                         �C@<���D�?            �@@       �                       @3�@��s����?             5@       �                         �B@����X�?             ,@       �                          A@      �?              @       �                          �@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     A@              &                    �?(*B���?E            @]@                                �?�+$�jP�?B             [@       	      
                   !@����e��?*            �P@        ������������������������       �                     �?        ������������������������       �        )            @P@                                 �?��6���?             E@                               �8@J�8���?             =@        ������������������������       �                     @                                �G@R�}e�.�?             :@                               �E@և���X�?
             ,@                               �B@z�G�z�?             $@                             ��v@�q�q�?             @                             �|Y<@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 �?�8��8��?             (@       ������������������������       �                     "@                              ���W@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @              %                   �?�	j*D�?             *@             $                  �E@X�<ݚ�?             "@              #                �̾w@և���X�?             @       !      "                  �4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        '      (                p�O@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M)KK��h2h3h4hVh<�h=Kub������������H�1�N�?oݟ�Kb�?R�Ω��?\��c�x�?�~�X��?��N̓�?xxxxxx�?�?UUUUUU�?UUUUUU�?              �?�������?333333�?              �?      �?        �9�s��?�c�1��?*.�u��?XG��).�?�������?333333�?      �?        ;�;��?vb'vb'�?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ���7���?Y�B��?      �?      �?      �?                      �?��y��y�?�a�a�?      �?        =��<���?�a�a�?<<<<<<�?�?      �?        �������?UUUUUU�?      �?      �?�������?�������?�������?UUUUUU�?      �?        �������?�������?      �?              �?              �?        �1���?*g���?l�l��?��I��I�?              �?;�;��?O��N���?�������?�������?�q�q�?�q�q�?              �?      �?                      �?              �?S��Ԧ6�?Y�JV���?�������?�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        E�pR���?u_[4�?��S�r
�??4և���?              �?�-��-��?�A�A�?�������?�������?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?vb'vb'�?;�;��?�<��<��?�a�a�?�q�q�?r�q��?      �?      �?      �?        ;�;��?ى�؉��?      �?      �?      �?      �?�m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?      �?              �?              �?      �?              �?                      �?      �?                      �?      �?        ���>4��?����S�?蝺���?���4>�?��18��?>�cp>�?d!Y�B�?ӛ���7�?              �?�?<<<<<<�?      �?      �?      �?                      �?      �?        #h8����?��c+���?              �?&���^B�?�%���^�?}g���Q�?AL� &W�?�ڕ�]��?��+Q��?�8��8��?9��8���?333333�?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?Y�B��?zӛ����?      �?      �?              �?�������?�������?      �?              �?      �?      �?        �������?�������?F]t�E�?/�袋.�?�������?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�z�G��?{�G�z�?ffffff�?�������?�������?�������?              �?      �?              �?        �������?333333�?      �?              �?      �?              �?      �?        �%N���?Ai�
��?�������?�������?>���>�?|���?wwwwww�?�?I�$I�$�?۶m۶m�?R���Q�?���Q��?�������?�������?      �?      �?      �?                      �?              �?�������?�������?      �?        �������?UUUUUU�?9��8���?�q�q�?      �?      �?      �?        �m۶m��?�$I�$I�?      �?              �?              �?                      �?      �?        �$I�$I�?�m۶m��?      �?                      �?�[���?d �?�*�?�������?�?UUUUUU�?UUUUUU�?      �?        �������?333333�?              �?      �?              �?      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ��P^Cy�?^Cy�5�?      �?        ------�?�������?<<<<<<�?�?�s�9��?�c�1Ƹ?      �?        ��Moz��?Y�B��?      �?      �?              �?�������?�?;�;��?;�;��?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        ]]]]]]�?�?              �?�>Q=h��?3	v�ܰ?�՝VwZ�?�RKE,�?UUUUUU�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?�Mozӛ�?d!Y�B�?UUUUUU�?UUUUUU�?      �?        ��8��8�?�q�q�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        �E]t��?t�E]t�?�������?�������?      �?      �?      �?        ��[��[�?�A�A�?      �?        �؉�؉�?;�;��?              �?���Q��?{�G�z�?�������?�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        ��L���?L�Ϻ��?      �?      �?      �?                      �?|���?|���?z��y���?�a�a�?�m۶m��?�$I�$I�?      �?      �?      �?      �?              �?      �?              �?              �?      �?      �?              �?              �?        ��Y��Y�?��)��)�?B{	�%��?/�����?|���?�>����?      �?                      �?=��<���?b�a��?|a���?�rO#,��?      �?        �;�;�?'vb'vb�?۶m۶m�?�$I�$I�?�������?�������?UUUUUU�?UUUUUU�?�������?333333�?              �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?vb'vb'�?;�;��?r�q��?�q�q�?۶m۶m�?�$I�$I�?      �?      �?              �?      �?                      �?      �?              �?        r�q��?�q�q�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�%\hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������       X                    �?�,�٧��?�           8�@               %                     @~��|��?�            pq@                                   �?l{��b��?W            �c@              	                    �?ДXࣿ?I             a@                                03�=@���7�?             F@                                �I5@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �A@        
                          @K@�c:��?/             W@                                  :@���L��?.            �V@                                  �B@�MI8d�?            �B@                                  �?ףp=
�?             >@                                 �7@H%u��?             9@                                  <@r�q��?             2@                                  �6@և���X�?             @        ������������������������       �                     @                                  �'@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     @                                  @F@և���X�?             @                                 �3@      �?             @        ������������������������       �                      @                                  �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     K@        ������������������������       �                     �?        !       $                     �?��2(&�?             6@        "       #                    $@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        &       W                   @B@b�
�p��?M            @^@       '       (                    @�q�QQ�?F            @[@        ������������������������       �                     *@        )       *                    )@     ��?>             X@        ������������������������       �                     @        +       <                    �?�?a/���?9            @V@        ,       9                    �?$G$n��?            �B@        -       8                    @�θ�?	             *@       .       /                 �&�)@      �?             (@        ������������������������       �                     @        0       7                  S�2@�q�q�?             "@       1       4                 ���,@և���X�?             @        2       3                   �-@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        5       6                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        :       ;                 ���@�8��8��?             8@        ������������������������       �                      @        ������������������������       �                     6@        =       V                 ���5@
j*D>�?              J@       >       O                 �|�<@D^��#��?            �D@       ?       J                 P�@��S���?             >@        @       C                   �2@r�q��?             (@        A       B                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        D       E                 pf�@ףp=
�?             $@        ������������������������       �                     @        F       I                 �&B@r�q��?             @        G       H                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        K       N                 ��/@�<ݚ�?	             2@       L       M                    3@      �?             0@        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                      @        P       Q                 pf�$@���!pc�?	             &@        ������������������������       �                      @        R       S                 03�1@�����H�?             "@       ������������������������       �                     @        T       U                 03C3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     (@        Y       �                     �?�ӭ�a��?            {@        Z       m                    �?VP��g��?5             W@        [       \                 ��";@j���� �?             A@        ������������������������       �                      @        ]       l                   �H@      �?             @@       ^       k                 X�l@@
;&����?             7@       _       j                    :@ҳ�wY;�?             1@       `       a                 Ȉ�P@���Q��?             $@        ������������������������       �                      @        b       i                    �?      �?              @       c       h                    �?�q�q�?             @       d       e                 0�HU@���Q��?             @        ������������������������       �                      @        f       g                 �U�X@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        n       o                    0@^l��[B�?!             M@        ������������������������       �                      @        p       q                 ��$:@����>4�?             L@        ������������������������       �                     "@        r       s                 03k:@��|�5��?            �G@        ������������������������       �                      @        t       �                    �?z�G�z�?            �F@       u       v                 �|Y>@���"͏�?            �B@        ������������������������       �                     $@        w       ~                   �E@�q�q�?             ;@        x       {                   @B@և���X�?             @        y       z                 0��J@      �?             @        ������������������������       �                      @        ������������������������       �                      @        |       }                  x#J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               �                   @H@      �?             4@        �       �                   �F@�C��2(�?             &@        �       �                 ���K@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���T@X�<ݚ�?             "@       �       �                 `fF<@����X�?             @       �       �                   �J@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���@hS>)��?�            @u@        ������������������������       �                     >@        �       �                 ��@ 7/��'�?�            `s@        ������������������������       �                      @        �       �                    �?ި�?�            @s@       �       �                 0C�E@��O���?�            �o@       �       �                 `�X#@h�N?���?�            @o@       �       �                   @@@��C[���?l             e@       �       �                 ���"@���Q�?^            �b@       �       �                   �>@�Z��L��?Y            �a@       �       �                 �|Y=@pH����?T            �`@       �       �                    �?؇���X�?-            �Q@        ������������������������       �                     @        �       �                   �3@�C��2(�?+            �P@        �       �                   �1@��s����?             5@        �       �                   �0@؇���X�?             @       �       �                 pFD!@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@d}h���?	             ,@        ������������������������       �                     @        �       �                   �2@�q�q�?             "@        �       �                 ��Y @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 0S5 @���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                 pf� @`Ӹ����?            �F@       ������������������������       �                    �C@        �       �                   �:@�q�q�?             @        ������������������������       �                     @        �       �                    <@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?'             P@       �       �                    �?      �?             @@       �       �                 �|�=@$�q-�?             *@       �       �                 ���@�C��2(�?	             &@        ������������������������       �                     @        �       �                 p&�@؇���X�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             3@        �       �                  sW@     ��?             @@        �       �                 ��,@      �?              @        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     8@        �       �                   �?@      �?              @        �       �                 pff@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �<@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     3@        �       �                   �7@ 7���B�?8            @T@       �       �                     @P���Q�?+             N@       �       �                   �)@���N8�?             E@        ������������������������       �        
             0@        �       �                    �?$�q-�?             :@        ������������������������       �                     @        �       �                    @@ףp=
�?             4@        ������������������������       �                     "@        �       �                   �*@"pc�
�?
             &@       �       �                   �F@      �?              @       �       �                   �A@���Q��?             @        ������������������������       �      �?              @        �       �                   �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�X�<ݺ?             2@        �       �                 �|Y<@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     5@        �       �                 ��?P@���Q��?             @        �       �                 �|�>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    :@�c�����?!            �J@       �       �                    �?r�q��?             8@        ������������������������       �                     @        �       �                    #@�ՙ/�?             5@        ������������������������       �                      @        ������������������������       �                     *@        �       �                    @ 	��p�?             =@        �       �                 ��yE@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     9@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������&��jq�?:�g *�?Hy�G�?n��n�?�&��jq�?${�ґ�?������?�������?F]t�E�?�.�袋�?�q�q�?9��8���?              �?      �?                      �?8��Moz�?Y�B���?��?>��=���?L�Ϻ��?��L���?�������?�������?���Q��?)\���(�?UUUUUU�?�������?۶m۶m�?�$I�$I�?              �?      �?      �?              �?      �?                      �?              �?              �?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?              �?      �?                      �?              �?      �?        t�E]t�?��.���?t�E]t�?F]t�E�?      �?                      �?              �?3(&ޏ�?�k����?������?�:#s��?              �?      �?      �?      �?        ���d%+�?7��Mmj�?���L�?к����?�؉�؉�?ى�؉��?      �?      �?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?b'vb'v�?;�;��?�]�ڕ��?,Q��+�?�?�������?UUUUUU�?�������?      �?      �?              �?      �?        �������?�������?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?9��8���?�q�q�?      �?      �?              �?      �?                      �?t�E]t�?F]t�E�?      �?        �q�q�?�q�q�?              �?      �?      �?      �?                      �?      �?              �?        �q�q�?�8��8��?�Mozӛ�?-d!Y��?�������?ZZZZZZ�?              �?      �?      �?�Mozӛ�?Y�B��?�������?�������?�������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?                      �?      �?        �=�����?��=���?              �?n۶m۶�?I�$I�$�?      �?        br1���?x6�;��?              �?�������?�������?v�)�Y7�?*�Y7�"�?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?]t�E�?F]t�E�?�������?�������?UUUUUU�?UUUUUU�?      �?              �?        r�q��?�q�q�?�m۶m��?�$I�$I�?�������?�������?              �?      �?              �?      �?              �?      �?                      �?      �?        TTTTTT�?]]]]]]�?      �?        �K��d��?Цm�?              �?��g�'�?S{����?�������?�?�v��/�?�I+��?�wɃg�?�B���Ǽ?�%�X��?7�i�6�?���.�d�?��Vؼ?�1���?z�rv��?۶m۶m�?�$I�$I�?              �?]t�E�?F]t�E�?z��y���?�a�a�?۶m۶m�?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?        I�$I�$�?۶m۶m�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?        ?�>��?l�l��?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?�؉�؉�?;�;��?]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?              �?              �?              �?      �?      �?      �?      �?              �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?              �?      �?      �?                      �?      �?        	�%����?h/�����?ffffff�?�������?��y��y�?�a�a�?      �?        �؉�؉�?;�;��?      �?        �������?�������?      �?        /�袋.�?F]t�E�?      �?      �?333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?        ��8��8�?�q�q�?۶m۶m�?�$I�$I�?      �?                      �?      �?              �?        333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �V�9�&�?:�&oe�?UUUUUU�?UUUUUU�?              �?�<��<��?�a�a�?              �?      �?        ������?�{a���?      �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ2�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                  x#J@"��p�?�           8�@                                  @��n:���?w           ��@                                    @�d�����?             C@        ������������������������       �                     3@               
                    �?�\��N��?             3@                                   @      �?              @        ������������������������       �                     @               	                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   @"pc�
�?             &@                                  �?ףp=
�?             $@        ������������������������       �                      @                                   �?      �?              @                                  @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               o                     @|����m�?`           `�@               .                 �|Y=@�&]�t��?�            �j@               #                    �?�r*e���?,            �R@                               ��*@�8��8��?             H@                                `f�)@�z�G��?             $@       ������������������������       �                     @                                   :@      �?             @                                  5@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                    :@P�Lt�<�?             C@       ������������������������       �                     ?@        !       "                   �6@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        $       )                    :@ȵHPS!�?             :@       %       (                    4@��S�ۿ?
             .@        &       '                   �2@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        *       -                   �;@"pc�
�?             &@        +       ,                   @<@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        /       n                    @��i]��?W            �a@       0       C                    �?�g+�v�?V             a@        1       2                    �?ףp=
�?             >@        ������������������������       �                      @        3       B                    �? �Cc}�?             <@       4       7                   �'@�LQ�1	�?             7@        5       6                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        8       9                     �?�����?             5@        ������������������������       �                     @        :       ;                   @B@�r����?             .@        ������������������������       �                      @        <       =                   �*@����X�?             @        ������������������������       �                     �?        >       ?                    5@r�q��?             @       ������������������������       �                     @        @       A                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        D       m                   @R@�NW���?@            �Z@       E       l                    �?��S�ۿ??            @Z@       F       G                   �)@���F6��?:            �X@        ������������������������       �                     7@        H       O                    �?@݈g>h�?.             S@        I       J                 ���<@@4և���?             ,@        ������������������������       �                     @        K       N                 ���=@      �?              @        L       M                 X��E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        P       [                   �*@��a�n`�?&             O@        Q       R                 �|�=@      �?              @        ������������������������       �                     �?        S       V                   @B@����X�?             @        T       U                    @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        W       X                   @D@z�G�z�?             @        ������������������������       �                      @        Y       Z                   �F@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        \       ]                 `fF:@�X�<ݺ?             K@        ������������������������       �        
             8@        ^       k                   �>@ףp=
�?             >@        _       j                   �<@�θ�?
             *@       `       i                     �?r�q��?	             (@       a       h                   �J@"pc�
�?             &@        b       c                 �|�?@���Q��?             @        ������������������������       �                      @        d       e                   �C@�q�q�?             @        ������������������������       �                     �?        f       g                    H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        p       �                 ��Y7@�<ݚ�?�            `u@       q       �                    �?���h���?�            s@        r       �                    �?��H���?<            @Y@       s       �                 �|�=@D�]�+��?:            �X@       t       �                    �?R�����?1             T@        u       �                    �?�Q����?             D@       v       y                    �?�ʻ����?             A@        w       x                 �&�)@      �?              @        ������������������������       �                     @        ������������������������       �                     @        z       �                 �&�)@�n_Y�K�?             :@       {       �                   �7@\X��t�?             7@        |                           5@؇���X�?             @       }       ~                 �{@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 ���@      �?             0@        ������������������������       �                     @        �       �                 ��� @���Q��?             $@       �       �                   @@X�<ݚ�?             "@        �       �                 �|=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �|Y=@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��g2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?���Q��?             D@        �       �                 ���@���7�?             6@        ������������������������       �                     �?        ������������������������       �                     5@        �       �                 �|Y=@r�q��?             2@        �       �                    ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   `3@�r����?             .@       ������������������������       �        
             *@        ������������������������       �                      @        ������������������������       �        	             2@        ������������������������       �                     @        �       �                 �|�=@��hJ,�?�            �i@       �       �                  s@�1�hP	�?d            �a@        ������������������������       �                     6@        �       �                    �?�8'��?U            @^@       �       �                    )@POͳF��?S            �]@        �       �                 ��|2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��-�=��?Q            @]@        �       �                   �4@�LQ�1	�?             7@        �       �                    3@؇���X�?             @       �       �                 `F�+@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?     ��?             0@       �       �                   �@      �?             ,@        �       �                 ���@r�q��?             @        ������������������������       �                     @        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        �       �                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �)@      �?              @       �       �                   �8@؇���X�?             @        ������������������������       �                     @        �       �                    ;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �4@`�q�0ܴ?@            �W@        �       �                 ��Y @@4և���?             <@       �       �                 P�@�r����?             .@       ������������������������       �                     $@        �       �                 @3�@���Q��?             @        ������������������������       �      �?              @        �       �                   �1@�q�q�?             @        ������������������������       �                     �?        �       �                   �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             *@        �       �                 �?$@Pa�	�?+            �P@        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                 pf�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �<@ ������?(            �O@        ������������������������       �                     @@        �       �                 ���"@�g�y��?             ?@       ������������������������       �                     :@        �       �                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�jTM��?&            �N@       �       �                 �&B@�BbΊ�?$             M@        ������������������������       �                     2@        �       �                    �?      �?             D@        �       �                 03�1@      �?              @       �       �                 `f�/@����X�?             @       �       �                    A@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �@     ��?             @@        ������������������������       �                     @        �       �                   �?@>���Rp�?             =@        �       �                 �?�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 @3�@�LQ�1	�?             7@        �       �                   @C@      �?             (@       ������������������������       �                     @        �       �                 �?�@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                    �B@        �                       `fmj@��Sݭg�?M            @]@       �       �                    �?�����?C            �X@       �       �                 ���Q@`Jj��?+             O@        �       �                 @3[Q@��s����?             5@       ������������������������       �        
             1@        ������������������������       �                     @        ������������������������       �                    �D@        �                           �?X�<ݚ�?             B@       �                         @I@�q�q�?             >@       �                       ���a@������?             ;@       �                          �?�θ�?             :@       �       �                   �8@����X�?             5@        ������������������������       �                      @        �                       `f^@���y4F�?             3@       �       
                p"�X@      �?
             0@                              0�"K@z�G�z�?	             .@                                 @@�q�q�?             @        ������������������������       �                      @                              `�iJ@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                �D@�����H�?             "@       ������������������������       �                     @              	                ЈT@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 �?�\��N��?
             3@        ������������������������       �                     "@        ������������������������       �                     $@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������J54v��?l�����?R�Ω��?\��c�x�?y�5���?Cy�5��?              �?y�5���?�5��P�?      �?      �?              �?      �?      �?      �?                      �?/�袋.�?F]t�E�?�������?�������?      �?              �?      �?�������?�������?      �?                      �?      �?                      �?�1O��?���a���?�+J�#�?�ީk9��?�u�)�Y�?0E>�S�?UUUUUU�?UUUUUU�?333333�?ffffff�?              �?      �?      �?      �?      �?              �?      �?                      �?(�����?���k(�?              �?�$I�$I�?۶m۶m�?      �?                      �?��N��N�?�؉�؉�?�������?�?�������?UUUUUU�?      �?                      �?      �?        /�袋.�?F]t�E�?�m۶m��?�$I�$I�?      �?                      �?      �?        _�_��?B�A��?�������?xxxxxx�?�������?�������?              �?۶m۶m�?%I�$I��?Y�B��?��Moz��?      �?      �?              �?      �?        �a�a�?=��<���?              �?�?�������?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?萚`���?�x+�R�?�������?�?�v�ļ�?ogH���?      �?        �P^Cy�?Cy�5��?n۶m۶�?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �s�9��?�c�1Ƹ?      �?      �?              �?�m۶m��?�$I�$I�?      �?      �?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        ��8��8�?�q�q�?      �?        �������?�������?ى�؉��?�؉�؉�?�������?UUUUUU�?/�袋.�?F]t�E�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?                      �?      �?              �?                      �?              �?9��8���?�q�q�?$����?pk�$��?T� w�l�?Y�&�?}h����?/����?�������?333333�?�������?ffffff�?�������?<<<<<<�?      �?      �?              �?      �?        ;�;��?ى�؉��?!Y�B�?��Moz��?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?      �?      �?      �?        333333�?�������?r�q��?�q�q�?      �?      �?      �?                      �?333333�?�������?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?F]t�E�?�.�袋�?      �?                      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?�������?�?      �?                      �?      �?                      �?KKKKKK�?�������?��^���?x��gں?      �?        N�zv�?�eP*L��?]�\��?e�e��?      �?      �?              �?      �?        }˷|˷�?�A�A�?Nozӛ��?d!Y�B�?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?              �?      �?      �?      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ��F}g��?W�+�ɥ?n۶m۶�?�$I�$I�?�������?�?      �?        333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        |���?|���?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?��}��}�?AA�?      �?        ��{���?�B!��?      �?        �������?�������?              �?      �?                      �?�y��!�?.�u�y�?�{a��?���=��?      �?              �?      �?      �?      �?�$I�$I�?�m۶m��?�������?333333�?              �?      �?                      �?      �?              �?      �?              �?�i��F�?GX�i���?UUUUUU�?UUUUUU�?      �?                      �?��Moz��?Y�B��?      �?      �?      �?        �������?333333�?      �?                      �?      �?              �?              �?        �i�i�?�|˷|��?����X�?^N��)x�?�B!��?���{��?�a�a�?z��y���?              �?      �?                      �?�q�q�?r�q��?UUUUUU�?UUUUUU�?{	�%���?B{	�%��?�؉�؉�?ى�؉��?�$I�$I�?�m۶m��?      �?        (������?6��P^C�?      �?      �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �q�q�?�q�q�?              �?      �?      �?              �?      �?              �?                      �?              �?      �?              �?              �?        y�5���?�5��P�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��(.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       T                    �?e�L��?�           8�@               !                    �?�,����?|            �h@                                    @$�3c�s�?8            �W@                                   �? qP��B�?            �E@              
                    �?(;L]n�?             >@                                 �H@ �q�q�?             8@       ������������������������       �                     3@               	                    J@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@                                   �?��x_F-�?            �I@                                  &@�ʈD��?            �E@                                  �@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                                ���@�}�+r��?             C@                                �|Y5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?������?             B@                                ���,@؇���X�?             @        ������������������������       �                     @                                P�h2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     =@                                    �?      �?              @                                �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        "       +                 03s@r�{o43�?D            �Y@        #       *                 ���@�7��?            �C@        $       )                    �?�r����?	             .@       %       &                 03S@8�Z$���?             *@        ������������������������       �                      @        '       (                   �7@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     8@        ,       1                 �y�'@     8�?+             P@        -       0                    �?�<ݚ�?             "@       .       /                 �|Y=@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        2       S                    I@^(��I�?&            �K@       3       4                 ��K.@p�v>��?             �G@        ������������������������       �                     @        5       6                 ��.@�q�q�?             E@        ������������������������       �                     @        7       R                   @F@�(�Tw��?            �C@       8       E                     �?���"͏�?            �B@        9       D                 `�&e@p�ݯ��?             3@       :       ?                 �|�;@      �?	             ,@        ;       >                   �5@؇���X�?             @        <       =                   �1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        @       A                   @@@؇���X�?             @        ������������������������       �                     @        B       C                   �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        F       Q                 03�7@�����H�?             2@        G       L                    �?      �?              @        H       I                    /@z�G�z�?             @        ������������������������       �                      @        J       K                 �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        M       P                    �?�q�q�?             @       N       O                   `3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        U       �                     @��*���?G           �@        V       W                   �1@vN#��?�            �j@        ������������������������       �                     1@        X       k                    �?@���S��?�            �h@        Y       Z                     �?p��@���?4            @U@        ������������������������       �                     ?@        [       j                    6@�����H�?"             K@       \       i                   @4@V�a�� �?             =@       ]       f                   �B@ȵHPS!�?             :@       ^       _                 `f�)@�X�<ݺ?             2@        ������������������������       �                     @        `       e                    :@�8��8��?	             (@        a       b                    5@      �?             @        ������������������������       �                      @        c       d                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        g       h                   �C@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     9@        l       �                     �?�X�C�?P             \@        m       �                   �R@�����?$            �H@       n       �                    �?t/*�?#            �G@       o       r                   �<@��s����?              E@        p       q                 `f�D@      �?             @        ������������������������       �                      @        ������������������������       �                      @        s       x                   @@@�S����?             C@        t       w                   �>@�}�+r��?             3@        u       v                   @>@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             (@        y       �                 03�U@�d�����?             3@       z                          @A@@�0�!��?             1@       {       |                 `fF:@      �?              @        ������������������������       �                     @        }       ~                   @M@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @A@���N8�?,            �O@       �       �                    �?$�q-�?            �C@       �       �                    1@�#-���?            �A@       �       �                   �@@ܷ��?��?             =@       �       �                    4@�>����?             ;@        �       �                    &@      �?              @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 �|Y=@�}�+r��?             3@       ������������������������       �        	             &@        �       �                 �|Y>@      �?              @       �       �                    @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     8@        �       �                    �?���I��?�            �r@        �       �                    �?������?0            @U@       �       �                   �>@N1���?!            �N@       �       �                    @����3��?             J@        ������������������������       �                     @        �       �                   �@���j��?             G@        �       �                 �&B@�n_Y�K�?             *@       �       �                 pf�@      �?              @        �       �                 �|Y:@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    3@6YE�t�?            �@@        �       �                 `f&+@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �:@ �Cc}�?             <@        ������������������������       �                     (@        �       �                   �;@     ��?
             0@        ������������������������       �                     �?        �       �                 �|�=@�r����?	             .@       �       �                    �?�8��8��?             (@        �       �                 �|�<@r�q��?             @        ������������������������       �                     �?        �       �                 pf&(@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   P2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    @r�q��?             8@       �       �                 �̼6@���y4F�?             3@        ������������������������       �                      @        �       �                 ��p@@�t����?	             1@        �       �                    @      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �       �                   �0@��6G���?�            �j@        �       �                 03�0@�eP*L��?             6@        ������������������������       �                     @        �       �                    �?z�G�z�?
             .@        ������������������������       �                     @        �       �                 ��<8@�q�q�?             "@        ������������������������       �                     �?        �       �                    @      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �?�@�0p<���?y             h@        �       �                 �Yu@��4+̰�?<            @X@       �       �                    7@�8���?&             M@        ������������������������       �                     8@        �       �                 ��L@l��\��?             A@       �       �                   �8@      �?             @@        �       �                 �&b@z�G�z�?             @        ������������������������       �                     @        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 X�l@@ 7���B�?             ;@       �       �                 ���@@4և���?
             ,@       ������������������������       �                      @        �       �                 �|�<@r�q��?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     *@        �       �                    >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �C@        �       �                 @3�@�8��8��?=             X@        �       �                    :@����X�?             @        ������������������������       �                      @        �       �                   �?@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        �       �                    (@���M�?7            @V@       �       �                 @Q!@�j��b�?$            �M@       �       �                 ��i @l��\��?             A@       �       �                   �3@ףp=
�?             >@        ������������������������       �                     @        ������������������������       �                     ;@        ������������������������       �                     @        �       �                   �:@H%u��?             9@        ������������������������       �                     (@        �       �                   �;@�θ�?             *@        ������������������������       �                      @        �       �                 �|�=@�C��2(�?             &@       ������������������������       �                      @        �       �                    A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     >@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������v�S(��?��X��?q�)`>��?G5���7�?x6�;��?1���\A�?�}A_З?��}A�?�?�������?UUUUUU�?�������?              �?�������?�������?      �?                      �?              �?              �?�?�������?�}A_з?A_���?�������?333333�?              �?      �?        (�����?�5��P�?      �?      �?              �?      �?        �q�q�?�q�q�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?      �?              �?      �?              �?        C����?���O ��?��[��[�?�A�A�?�������?�?;�;��?;�;��?      �?        /�袋.�?F]t�E�?              �?      �?              �?              �?             ��?      �?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?�7�}���?J��yJ�?ڨ�l�w�?L� &W�?      �?        UUUUUU�?UUUUUU�?              �?�o��o��?� � �?v�)�Y7�?*�Y7�"�?^Cy�5�?Cy�5��?      �?      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �q�q�?�q�q�?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?      �?        ����?�+�+�+�?z����f�?C�(��L�?              �?���^K�?/,FBi��?�?�������?              �?�q�q�?�q�q�?a���{�?��{a�?�؉�؉�?��N��N�?�q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?      �?                      �?�$I�$I�?n۶m۶�?^N��)x�?����X�?�;����?W�+���?z��y���?�a�a�?      �?      �?              �?      �?        (������?^Cy�5�?�5��P�?(�����?۶m۶m�?�$I�$I�?      �?                      �?      �?        Cy�5��?y�5���?ZZZZZZ�?�������?      �?      �?      �?        �������?333333�?              �?      �?              �?                      �?      �?                      �?��y��y�?�a�a�?�؉�؉�?;�;��?�A�A�?_�_�?��=���?a���{�?�Kh/��?h/�����?      �?      �?      �?      �?      �?        �5��P�?(�����?      �?              �?      �?�������?�������?      �?                      �?      �?              �?      �?      �?              �?              �?        Y�%�X�?�6�i��?�������?�?�:ڼO�?�}�K�`�?��N��N�?'vb'vb�?              �?ozӛ���?!Y�B�?ى�؉��?;�;��?      �?      �?      �?      �?              �?      �?              �?                      �?'�l��&�?e�M6�d�?333333�?�������?              �?      �?        %I�$I��?۶m۶m�?      �?              �?      �?              �?�������?�?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?        �������?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?UUUUUU�?6��P^C�?(������?              �?<<<<<<�?�?      �?      �?              �?      �?              �?              �?        �������?��0�?t�E]t�?]t�E�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        ��3-�?�O�l.�?_\����? tT����?j��FX�?a���{�?      �?        ------�?�������?      �?      �?�������?�������?      �?              �?      �?              �?      �?        	�%����?h/�����?n۶m۶�?�$I�$I�?      �?        �������?UUUUUU�?      �?              �?      �?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?      �?��^����?�E(B�?�N��?��/���?------�?�������?�������?�������?              �?      �?              �?        )\���(�?���Q��?      �?        ى�؉��?�؉�؉�?              �?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJx�+hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       P                    �?��ϙLq�?�           8�@                                   �?��g�ao�?^            �a@                                0Cd=@�y��*�?'             M@                                P��+@�X����?             6@        ������������������������       �                     @                                �|Y=@��S���?	             .@                                 �-@�z�G��?             $@        ������������������������       �                      @        	       
                     @      �?              @        ������������������������       �                     �?                                  �0@؇���X�?             @        ������������������������       �                     @                                03�-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 S�2@z�G�z�?             @        ������������������������       �                      @                                ��9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     B@               %                   �:@ҳ�wY;�?7            @U@               $                    �?8����?             7@                                  3@�q�q�?             5@                                �	N@���Q��?             @                               ��}@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @               !                   @7@      �?
             0@                                 ��y@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        "       #                 xF*@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        &       ?                     �?��a�n`�?(             O@        '       >                    �?f���M�?             ?@       (       =                    I@
j*D>�?             :@       )       :                    �?�G��l��?             5@       *       5                  xCH@     ��?             0@       +       2                   @@@      �?              @       ,       1                 �|�=@r�q��?             @       -       .                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        /       0                 ��2>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        3       4                   �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        6       7                 0�c@      �?              @       ������������������������       �                     @        8       9                 X�,@@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ;       <                 �;�p@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        @       C                 �|Y=@��a�n`�?             ?@        A       B                 ��Y&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        D       E                     @ 	��p�?             =@        ������������������������       �                     @        F       O                 �|Y?@HP�s��?             9@       G       L                  S�'@�����H�?             2@       H       I                 ���@      �?	             0@        ������������������������       �                      @        J       K                   @@      �?              @       ������������������������       �z�G�z�?             @        ������������������������       �                     @        M       N                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        Q       �                    �?V��	3�?g           ��@        R       �                 �D�H@�$�q��?n             e@       S       f                     @ XөM"�?Y             a@        T       U                     �?h�WH��?"             K@        ������������������������       �                     @        V       W                 `f�)@`�H�/��?             �I@        ������������������������       �        
             0@        X       e                    :@؇���X�?            �A@       Y       ^                   �3@�GN�z�?             6@       Z       ]                   �*@�C��2(�?	             &@       [       \                    <@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        _       d                    D@���|���?             &@       `       c                    �?      �?              @       a       b                    <@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     *@        g       z                  SE"@��q7L��?7            �T@        h       w                    �?��R[s�?            �A@       i       j                    8@     ��?             @@        ������������������������       �                     *@        k       l                 ���@p�ݯ��?             3@        ������������������������       �                      @        m       t                 �̌@�t����?             1@       n       o                 ��@�C��2(�?	             &@       ������������������������       �                     @        p       q                    �?      �?             @        ������������������������       �                      @        r       s                   �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        u       v                 ��� @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        x       y                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        {       �                 ���1@�q�q�?             H@        |       }                   �&@��.k���?             1@        ������������������������       �                     @        ~       �                    �?z�G�z�?	             $@              �                   �D@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�n`���?             ?@        ������������������������       �                     &@        �       �                 �̼6@�z�G��?             4@        ������������������������       �                      @        �       �                 ��T?@�<ݚ�?             2@       ������������������������       �                     &@        �       �                    %@և���X�?             @        ������������������������       �                     @        �       �                 pf�C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    !@     ��?             @@        ������������������������       �                     �?        �       �                  DpR@`Jj��?             ?@        �       �                 ��\O@؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     1@        �       �                 `f^4@Ԫ2��?�            �x@       �       �                    �?$�q-�?�            q@       �       �                    �?��u���?�            pp@        �       �                 �|Y=@�>����?             ;@        �       �                  ��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        �       �                 0SE @�JM-Xy�?�            �m@       �       �                   @4@@v�禺�?T            �`@        �       �                   �2@d}h���?             ,@        ������������������������       �                     @        �       �                   �3@���!pc�?	             &@        �       �                 �?�@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        �       �                 P�@r�q��?             @       ������������������������       �                     @        �       �                 @3�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��) @�U�:��?H            �]@       �       �                 �?�@ 	��p�?G             ]@       �       �                 �?$@��
���?2            �R@       �       �                 ���@������?            �D@        ������������������������       �                     6@        �       �                    7@�KM�]�?             3@        ������������������������       �                     @        �       �                    9@؇���X�?             ,@        �       �                 `fF@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 pf�@�8��8��?	             (@       ������������������������       �                     @        �       �                 �|Y>@z�G�z�?             @       �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     A@        �       �                 @3�@�p ��?            �D@        �       �                    :@      �?             0@        ������������������������       �                     @        �       �                   �?@��
ц��?             *@        ������������������������       �                      @        �       �                   �A@���|���?             &@        ������������������������       �      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     9@        ������������������������       �                      @        �       �                   �3@ pƵHP�?<             Z@        �       �                   �2@���}<S�?             7@       ������������������������       �                     $@        �       �                     @8�Z$���?             *@        �       �                   �'@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �        .            @T@        �       �                    �?���Q��?             $@        ������������������������       �                     �?        �       �                    �?X�<ݚ�?             "@       �       �                    +@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    @�E��ӭ�?O            �_@        �       �                 ��T?@p�ݯ��?             3@       �       �                    �?�eP*L��?             &@       �       �                     @X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                 ���9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @      �?              @       ������������������������       �                     @        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                           �?�Ы܋��?C            �Z@       �                          �?���|���?#            �K@       �       �                    �?䯦s#�?!            �J@        ������������������������       �                     �?        �                          �>@�n_Y�K�?              J@        �       �                   �<@l��[B��?             =@        ������������������������       �                     @        �       �                 ��$:@��
ц��?             :@        ������������������������       �                     @        �       �                 03k:@�eP*L��?             6@        ������������������������       �                     @        �       �                 `fF<@�\��N��?             3@       �       �                 �|�?@���!pc�?             &@        ������������������������       �                     @        �       �                   �C@      �?              @        ������������������������       �                      @        �       �                    H@r�q��?             @        ������������������������       �                     @        �       �                   �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @>@      �?              @       �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                �;@��<b���?             7@                                 7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @              
                  @H@R���Q�?             4@                             03�U@��S�ۿ?             .@       ������������������������       �        	             *@              	                �w|c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              ���W@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                              �̌4@0G���ջ?              J@        ������������������������       �                     �?                                 �?`'�J�?            �I@                              03�7@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                              �T�I@`���i��?             F@       ������������������������       �                    �A@                                 ;@�����H�?             "@                                  @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������Ӭ����?�X�>��?��3m���?�
fI9 �?GX�i��?�4�rO#�?]t�E]�?�E]t��?              �?�������?�?333333�?ffffff�?      �?              �?      �?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?8��Moz�?d!Y�B�?UUUUUU�?UUUUUU�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?�$I�$I�?۶m۶m�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�c�1��?�s�9��?��RJ)��?��Zk���?b'vb'v�?;�;��?��y��y�?1�0��?      �?      �?      �?      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?      �?              �?      �?              �?      �?              �?      �?      �?      �?                      �?333333�?�������?      �?                      �?      �?              �?        �s�9��?�c�1Ƹ?      �?      �?              �?      �?        ������?�{a���?      �?        q=
ףp�?{�G�z�?�q�q�?�q�q�?      �?      �?      �?              �?      �?�������?�������?      �?              �?      �?      �?                      �?      �?        O�o�z2�?as �
��?pƵHP�?����W�?�d�*al�?�͂j���?B{	�%��?��^B{	�?              �?�?�������?              �?�$I�$I�?۶m۶m�?]t�E�?�袋.��?F]t�E�?]t�E�?�$I�$I�?۶m۶m�?      �?                      �?              �?F]t�E�?]t�E]�?      �?      �?UUUUUU�?�������?      �?                      �?              �?      �?                      �?��\V��?��FS���?PuPu�?X|�W|��?      �?      �?              �?Cy�5��?^Cy�5�?      �?        �������?�������?F]t�E�?]t�E�?              �?      �?      �?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?�������?�?      �?        �������?�������?      �?      �?              �?      �?              �?      �?              �?      �?        �9�s��?�c�1��?      �?        ffffff�?333333�?              �?9��8���?�q�q�?      �?        ۶m۶m�?�$I�$I�?              �?      �?      �?              �?      �?              �?      �?      �?        �B!��?���{��?�$I�$I�?۶m۶m�?              �?      �?                      �?$���>��?p�}��?�؉�؉�?;�;��?J�y�z��?��2�*��?�Kh/��?h/�����?UUUUUU�?UUUUUU�?      �?                      �?      �?        lE�pR��?��}ylE�?�d�M6��?6�d�M6�?I�$I�$�?۶m۶m�?      �?        F]t�E�?t�E]t�?333333�?�������?      �?        UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?              �?      �?              �?      �?        �A�I�?�pR�屵?������?�{a���?&�X�%�?O贁N�?p>�cp�?������?      �?        �k(���?(�����?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?        Q��+Q�?��+Q��?      �?      �?      �?        �;�;�?�؉�؉�?              �?]t�E]�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?'vb'vb�?;�;��?ӛ���7�?d!Y�B�?      �?        ;�;��?;�;��?      �?      �?UUUUUU�?UUUUUU�?      �?              �?              �?        333333�?�������?      �?        r�q��?�q�q�?۶m۶m�?�$I�$I�?              �?      �?              �?        �q�q�?r�q��?Cy�5��?^Cy�5�?t�E]t�?]t�E�?r�q��?�q�q�?              �?      �?              �?      �?              �?      �?              �?      �?              �?      �?      �?      �?                      �?��XQ�?蝺���?]t�E]�?F]t�E�?�����?�V�9�&�?      �?        ;�;��?ى�؉��?GX�i���?���=��?              �?�;�;�?�؉�؉�?      �?        ]t�E�?t�E]t�?              �?y�5���?�5��P�?F]t�E�?t�E]t�?      �?              �?      �?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?��,d!�?��Moz��?UUUUUU�?UUUUUU�?      �?                      �?333333�?333333�?�������?�?      �?              �?      �?              �?      �?        333333�?�������?      �?                      �?      �?        vb'vb'�?�؉�؉�?              �?�������?�?۶m۶m�?�$I�$I�?              �?      �?        F]t�E�?F]t�E�?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJH�SshG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������       
                    @�3)0�F�?�           8�@                                    @x�����?            �C@        ������������������������       �                     2@                                ��*4@�ՙ/�?             5@        ������������������������       �                     $@                                   �?���!pc�?             &@        ������������������������       �                     @               	                    @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @               �                   �R@�D���~�?�            �@              U                    �?\>��?�           ��@               D                    �?&� �N�?g             d@              /                 �|Y=@"Ae���?=            �W@               *                 0C�<@h+�v:�?             A@                                 P,@�q�����?             9@                                  @@���!pc�?	             &@                                ���@���Q��?             @        ������������������������       �                     �?                                   �?      �?             @        ������������������������       �                     �?                                  �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                    @X�Cc�?	             ,@                                  �9@      �?             @        ������������������������       �                      @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                )                    <@���Q��?             $@       !       (                     @      �?              @       "       #                    (@؇���X�?             @        ������������������������       �                     @        $       '                    �?      �?             @       %       &                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        +       ,                    �?�����H�?             "@       ������������������������       �                     @        -       .                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        0       A                 м�J@���*�?#             N@       1       2                 �?�-@H�ՠ&��?             K@       ������������������������       �                     5@        3       :                 ��-7@�'�`d�?            �@@        4       7                    �?�n_Y�K�?             *@        5       6                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        8       9                 `fv2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ;       @                    �?ףp=
�?             4@       <       =                    B@�����H�?
             2@        ������������������������       �                     &@        >       ?                   �F@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        B       C                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        E       T                    �?Pa�.l�?*            �P@       F       G                 �|Y=@�m����?%            �M@        ������������������������       �                     @        H       I                    �?X�Emq�?!            �J@        ������������������������       �                     5@        J       S                 X��A@      �?             @@       K       P                   `3@��S�ۿ?             >@       L       M                 ���@ 7���B�?             ;@        ������������������������       �                     @        N       O                 ��(@P���Q�?             4@       ������������������������       �@4և���?	             ,@        ������������������������       �                     @        Q       R                 03�7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        V       ]                    +@6T^�P4�?             {@        W       \                    '@��S���?
             .@       X       Y                 ���4@��
ц��?	             *@        ������������������������       �                     @        Z       [                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ^       �                    �?��N�Т�?           0z@        _       �                 ���P@      �?F             \@       `       �                    @�Ы܋��?C            �Z@       a       v                 `f�$@���B���?A             Z@        b       c                   �1@8�A�0��?             6@        ������������������������       �                     @        d       q                   �"@�\��N��?             3@       e       l                   �4@X�Cc�?             ,@        f       k                    �?�q�q�?             @       g       h                 �&B@z�G�z�?             @        ������������������������       �                     @        i       j                 xF� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        m       p                   �9@      �?              @       n       o                 pff@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        r       s                 Ь�#@z�G�z�?             @        ������������������������       �                     @        t       u                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        w       �                     @��1��?1            �T@       x       �                   �*@0�,���?'            �P@        y       �                   �J@�����?             5@       z                           �?P���Q�?             4@       {       |                   �B@�}�+r��?             3@       ������������������������       �        	             0@        }       ~                    F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     G@        �       �                    @���Q��?
             .@       �       �                    �?��
ц��?	             *@       �       �                    �?�z�G��?             $@       �       �                   �0@և���X�?             @       �       �                 @3�/@      �?             @       �       �                 ��Y.@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 03�1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?T�s�6&�?�            0s@       �       �                 ��$:@LzP��?�            Pq@       �       �                 ��@��[B��?�             m@        ������������������������       �                    �D@        �       �                     �? �r�ɻ?�            �g@        ������������������������       �                     �?        �       �                 �|Y=@�+?�?�            �g@       �       �                 ���$@Pa�	�?D            �X@       �       �                   �3@�\=lf�?.            �P@        �       �                 0S5 @�}�+r��?             3@        �       �                   �1@      �?              @        ������������������������       �                     �?        �       �                 �?�@؇���X�?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     &@        ������������������������       �                      H@        �       �                    &@      �?             @@        �       �                    5@      �?              @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     8@        �       �                     @|)����?<            �V@        �       �                 �|�=@ �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        �       �                    ?@pH����?)            �P@       �       �                  sW@�X�<ݺ?             B@        ������������������������       ��q�q�?             @        ������������������������       �                    �@@        �       �                   @@@�חF�P�?             ?@        �       �                   �@�q�q�?             "@        ������������������������       �                     �?        �       �                 �?�@      �?              @        ������������������������       �                      @        �       �                 ��I @�q�q�?             @        ������������������������       �      �?             @        ������������������������       �                      @        �       �                   @C@�C��2(�?             6@       ������������������������       �                     (@        �       �                 @3�@z�G�z�?             $@        �       �                 �?�@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                     �?f.i��n�?!            �F@       �       �                 `f�;@��V#�?            �E@        �       �                 03k:@�q�q�?	             (@        ������������������������       �                     �?        �       �                   �J@���|���?             &@       �       �                   @G@      �?              @       �       �                   �C@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                  x#J@�n`���?             ?@       �       �                   �>@؇���X�?             5@        �       �                   `H@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �A@��S�ۿ?             .@        ������������������������       �                      @        �       �                 ��yC@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `�iJ@�z�G��?             $@        ������������������������       �                     �?        �       �                 03�M@�<ݚ�?             "@       �       �                    A@����X�?             @       �       �                 `f�K@�q�q�?             @       �       �                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     >@        �       �                    �?z���=��?/            @S@       ������������������������       �        !            �K@        �       �                   �B@8�A�0��?             6@       �       �                    �?�	j*D�?             *@       �       �                    �?�q�q�?             "@       �       �                   �8@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                  "&d@      �?             @        ������������������������       �                      @        �       �                 @��v@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������Rl���?�[�'��?�A�A�?��o��o�?              �?�a�a�?�<��<��?              �?F]t�E�?t�E]t�?      �?        �������?333333�?      �?                      �?��y��y�?�0�0�?�Hm�Hm�?�n%�n%�?���2��?�l<�?�?�w6�;�?W�+���?xxxxxx�?�������?���Q��?�p=
ף�?t�E]t�?F]t�E�?333333�?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?%I�$I��?�m۶m��?      �?      �?      �?              �?      �?              �?      �?        333333�?�������?      �?      �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?              �?      �?              �?                      �?              �?�q�q�?�q�q�?              �?      �?      �?              �?      �?        """"""�?wwwwww�?������?{	�%���?      �?        6�d�M6�?'�l��&�?;�;��?ى�؉��?�$I�$I�?۶m۶m�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�q�q�?�q�q�?      �?        �m۶m��?�$I�$I�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        ��~5&�?5&����?��}ylE�?�V'u�?              �?5�x+��?�}�	��?              �?      �?      �?�������?�?	�%����?h/�����?      �?        ffffff�?�������?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ;~��_�?�Ł�@�?�������?�?�;�;�?�؉�؉�?              �?      �?      �?              �?      �?                      �?\��+��?I��/��?      �?      �?蝺���?��XQ�?ى�؉��?��؉���?/�袋.�?颋.���?              �?�5��P�?y�5���?�m۶m��?%I�$I��?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?�������?�������?      �?              �?      �?              �?      �?        ,Q��+�?�+Q���?g��1��?Ez�rv�?�a�a�?=��<���?�������?ffffff�?(�����?�5��P�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?333333�?�������?�;�;�?�؉�؉�?ffffff�?333333�?�$I�$I�?۶m۶m�?      �?      �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?              �?              �?        ��[&�d�?]0"��ش?��Z��?��o+��?a���{�?�i��F�?      �?        �ќ5(�?o��2�|�?      �?        \���%�?Fڱa��?|���?|���?"=P9���?g��1��?�5��P�?(�����?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?      �?              �?              �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?        ��/��/�?h�h��?�������?UUUUUU�?              �?      �?        �1���?z�rv��?��8��8�?�q�q�?UUUUUU�?UUUUUU�?      �?        �Zk����?��RJ)��?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        ]t�E�?F]t�E�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?        �`�`�?�>�>��?eMYS֔�?6eMYS��?UUUUUU�?UUUUUU�?              �?F]t�E�?]t�E]�?      �?      �?      �?      �?              �?      �?      �?              �?      �?        �9�s��?�c�1��?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?�������?�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        ffffff�?333333�?              �?9��8���?�q�q�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?              �?              �?              �?        
qV~B��?�cj`��?              �?颋.���?/�袋.�?;�;��?vb'vb'�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�8�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       P                    �?�_%����?�           8�@                                    @������?�            �o@                                  �?XB���?_             b@                               ��*@ ;=֦��?O            �^@                                  �J@ףp=
�?             >@                                  �? 	��p�?             =@        ������������������������       �                     @                                  �9@$�q-�?             :@        	       
                   �6@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  �'@���N8�?             5@        ������������������������       �                     "@                                  �B@�8��8��?             (@       ������������������������       �                     "@                                   D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        <             W@                                   @���}<S�?             7@        ������������������������       �                      @        ������������������������       �                     5@               -                    �?      �?J            �[@               &                    �?     ��?             @@                                   �?�eP*L��?
             &@                                �&�)@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                P��+@      �?              @        ������������������������       �                      @                !                   �@�q�q�?             @        ������������������������       �                     �?        "       #                   �7@z�G�z�?             @        ������������������������       �                      @        $       %                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        '       ,                    �?؇���X�?             5@       (       )                 �|�6@ףp=
�?             4@        ������������������������       �                      @        *       +                 ���@�����H�?             2@        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     �?        .       G                    �?�e����?/            �S@       /       4                 P�@      �?              M@        0       3                 ��@�8��8��?             (@       1       2                    A@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        5       @                    �?�û��|�?             G@       6       ;                 ��&@�q�q�?             ;@       7       8                 �|Y>@�����H�?	             2@       ������������������������       �                     ,@        9       :                    A@      �?             @        ������������������������       �                      @        ������������������������       �                      @        <       ?                 ���1@�<ݚ�?             "@       =       >                   �D@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        A       F                 ���4@�\��N��?             3@       B       C                    7@"pc�
�?             &@        ������������������������       �                     @        D       E                 `fv1@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        H       I                    @R���Q�?             4@        ������������������������       �                      @        J       K                    4@�X�<ݺ?             2@       ������������������������       �                     $@        L       O                    @      �?              @       M       N                 �|�:@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        Q       t                 �?�@��L#@r�?           �|@        R       a                    �?�c!�^�?\            @b@        S       T                 ��y@��2(&�?             6@        ������������������������       �                     �?        U       ^                   @@؇���X�?             5@       V       W                   @9@�r����?             .@        ������������������������       �                     �?        X       Y                 ���@@4և���?             ,@        ������������������������       �                     @        Z       [                 �|=@؇���X�?             @        ������������������������       �                     @        \       ]                 �|�=@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        _       `                 �|Y=@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        b       s                 �?$@�g�y��?O             _@       c       d                     @H�!b	�?4            @T@        ������������������������       �                     (@        e       f                 ���@p��%���?,            @Q@        ������������������������       �                     5@        g       h                 ���@�8��8��?             H@        ������������������������       �                      @        i       l                    �?�nkK�?             G@        j       k                  ��@�C��2(�?             &@        ������������������������       �                     @        ������������������������       �؇���X�?             @        m       n                 ��@��?^�k�?            �A@       ������������������������       �                     8@        o       p                 �|Y9@�C��2(�?             &@        ������������������������       �                     @        q       r                 �|Y>@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                    �E@        u       �                    @�q!I�?�            `s@        v       w                     @�q�q�?             ;@        ������������������������       �                      @        x       �                    @�\��N��?             3@       y       z                 ��|2@���Q��?
             .@        ������������������������       �                     @        {       |                    �?ףp=
�?             $@       ������������������������       �                     @        }       ~                     @�q�q�?             @        ������������������������       �                     �?               �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     �?������?�            �q@        �       �                    �?�JY�8��?A             Y@        �       �                 8�VQ@p�ݯ��?             C@       �       �                    �?؇���X�?             5@       �       �                 �|�;@     ��?
             0@        ������������������������       �                     �?        �       �                 ��";@�r����?	             .@        ������������������������       �                     �?        �       �                  �>@@4և���?             ,@        ������������������������       �                      @        �       �                 p�i@@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?ҳ�wY;�?             1@       �       �                   �5@�q�q�?             (@        ������������������������       �                      @        �       �                 p"�X@z�G�z�?             $@       ������������������������       �                     @        �       �                   @E@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 tՌs@���Q��?             @       �       �                    �?      �?             @        ������������������������       �                     �?        �       �                 �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @@Z��Yo��?)             O@        �       �                    <@�n_Y�K�?             :@        ������������������������       �                     @        �       �                   @>@\X��t�?             7@       �       �                 �|�?@X�<ݚ�?             2@        ������������������������       �                     @        �       �                   �9@��S���?             .@        ������������������������       �                      @        �       �                   @=@�n_Y�K�?
             *@       �       �                 `f�;@�eP*L��?	             &@       �       �                   �K@���Q��?             $@       �       �                 03k:@؇���X�?             @        ������������������������       �                     �?        �       �                    H@r�q��?             @       �       �                   �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?tk~X��?             B@       �       �                  x#J@�������?             >@       �       �                 `f�D@��S�ۿ?             .@        �       �                 �|�<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                 03�M@���Q��?
             .@        �       �                    7@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03�U@z�G�z�?             $@        ������������������������       �                     @        �       �                  �6f@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �                         @E@hau��?p            �f@       �       �                    �?0��^�?e            �d@        �       �                 м;4@���!pc�?             6@       �       �                    '@      �?	             (@        ������������������������       �                      @        �       �                     @���Q��?             $@        ������������������������       �                      @        �       �                 03�-@      �?              @        �       �                    3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                 �|�=@<�&9�?W             b@       �       �                   �+@�$��y��?:            @X@       �       �                    $@�r����?&             N@       �       �                 0SE @�C��2(�?             F@       �       �                 ��) @��s����?             5@       �       �                 @3�@R���Q�?             4@        �       �                   �4@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                    3@�r����?
             .@        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     7@        �       �                 �|�<@      �?	             0@       �       �                    4@؇���X�?             ,@        �       �                   �2@���Q��?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     "@        ������������������������       �                      @        �       �                    �?�?�|�?            �B@       �       �                 0��D@ 7���B�?             ;@       ������������������������       �                     8@        �       �                 ��?P@�q�q�?             @       �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                 @3�@�q�q�?             H@        �       �                   �?@      �?             (@        ������������������������       �                     �?        �       �                   �A@���!pc�?             &@       ������������������������       ��q�q�?             @        ������������������������       �z�G�z�?             @        �       �                   �>@4?,R��?             B@        �       �                    $@      �?             @        �       �                 �̌!@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �                           @��S�ۿ?             >@        �                         �3@��S�ۿ?	             .@                              `fF)@      �?              @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     @                              �TE@��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        ������������������������       �                     0@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������z���� �?@Bx��?�?xxxxxx�?�{a���?GX�i���?XG��).�?�%C��6�?�������?�������?�{a���?������?              �?;�;��?�؉�؉�?�������?�������?              �?      �?        �a�a�?��y��y�?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?d!Y�B�?ӛ���7�?      �?                      �?      �?      �?      �?      �?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?�������?�������?              �?�q�q�?�q�q�?      �?                      �?      �?        �-��-��?�A�A�?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?      �?                      �?8��Moz�?��,d!�?UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?              �?      �?              �?      �?        �q�q�?9��8���?      �?      �?              �?      �?              �?        y�5���?�5��P�?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        333333�?333333�?              �?��8��8�?�q�q�?      �?              �?      �?�������?�������?              �?      �?              �?        �YLg1��?���b:��?t�Ν;w�?Ĉ#F��?��.���?t�E]t�?      �?        ۶m۶m�?�$I�$I�?�������?�?              �?n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?      �?        �������?UUUUUU�?              �?      �?        ��{���?�B!��?b�2�tk�?�����H�?      �?        �g��%�?ہ�v`��?      �?        UUUUUU�?UUUUUU�?              �?�Mozӛ�?d!Y�B�?]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?_�_��?�A�A�?      �?        ]t�E�?F]t�E�?      �?        �������?UUUUUU�?      �?      �?      �?              �?        T�Cu;T�?X�x�W�?UUUUUU�?UUUUUU�?              �?�5��P�?y�5���?333333�?�������?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�F6���?��&���?)\���(�?�G�z��?^Cy�5�?Cy�5��?۶m۶m�?�$I�$I�?      �?      �?              �?�������?�?              �?n۶m۶�?�$I�$I�?      �?        �������?UUUUUU�?              �?      �?              �?        �������?�������?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?              �?      �?        �������?333333�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?!�B!�?���{��?ى�؉��?;�;��?              �?��Moz��?!Y�B�?r�q��?�q�q�?      �?        �������?�?      �?        ى�؉��?;�;��?]t�E�?t�E]t�?�������?333333�?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?              �?r�q��?9��8���?�������?�������?�������?�?      �?      �?              �?      �?              �?        333333�?�������?�������?�������?      �?                      �?�������?�������?      �?        333333�?�������?              �?      �?              �?        ��o���?��Y@�H�?y�oq�?×b@:�?F]t�E�?t�E]t�?      �?      �?      �?        �������?333333�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        EɮM���?��DɮM�?����?W?���?�������?�?]t�E�?F]t�E�?z��y���?�a�a�?333333�?333333�?�������?�������?      �?      �?      �?        �������?�?              �?      �?                      �?      �?              �?      �?۶m۶m�?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?*�Y7�"�?к����?	�%����?h/�����?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?              �?        �������?�������?      �?      �?              �?t�E]t�?F]t�E�?UUUUUU�?UUUUUU�?�������?�������?�8��8��?r�q��?      �?      �?      �?      �?      �?                      �?      �?        �������?�?�������?�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJUehG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM)hjh))��}�(h,h/h0M)��h2h3h4hph<�h=Kub������       �                     @|��;;��?�           8�@               %                    �?)O���?�            @t@                                03[=@PX�V|�?W            `a@                                03;<@�C��2(�?%            �P@                                 �;@      �?$             P@                                   �?H%u��?             9@                                  )@�θ�?             *@        ������������������������       �                     @        	       
                   �5@�q�q�?             "@        ������������������������       �                     �?                                ���*@      �?              @        ������������������������       �                      @                                ��m1@r�q��?             @        ������������������������       �                     @                                  �9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@                                `f�)@ ���J��?            �C@        ������������������������       �                     1@                                   �?���7�?             6@        ������������������������       �                      @                                  �*@P���Q�?             4@                                  �B@r�q��?             @       ������������������������       �                     @                                   D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             ,@        ������������������������       �                      @                                  "�b@ �й���?2            @R@       ������������������������       �        &             M@        !       "                    �?��S�ۿ?             .@        ������������������������       �                     @        #       $                 03c@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        &       C                 ��D:@��!w�K�?v             g@        '       >                    ,@�8��8��?5             U@       (       )                    @�1�`jg�?#            �K@        ������������������������       �                      @        *       =                   �*@=QcG��?            �G@       +       ,                    �?Du9iH��?            �E@        ������������������������       �                     �?        -       <                    �?@4և���?             E@       .       3                   �(@��(\���?             D@        /       2                    &@      �?
             0@       0       1                   �5@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                      @        4       9                   �C@�8��8��?             8@       5       6                 �|Y<@���N8�?             5@        ������������������������       �                     (@        7       8                 �|�=@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        :       ;                   �F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ?       @                    �?\-��p�?             =@       ������������������������       �                     6@        A       B                    :@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        D       �                    @Fn�圴�?A            @Y@       E       f                    �?`�Q��?@             Y@        F       [                 pVAH@�e����?            �C@       G       Z                 0�&C@����X�?             5@       H       Y                    �?և���X�?             ,@       I       J                 ��";@�n_Y�K�?
             *@        ������������������������       �                     �?        K       L                   �;@�q�q�?	             (@        ������������������������       �                      @        M       X                     �?z�G�z�?             $@       N       U                  �>@�<ݚ�?             "@       O       T                    �?؇���X�?             @       P       S                 X�lE@r�q��?             @        Q       R                 ��2>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        V       W                   �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        \       ]                 �|Y<@X�<ݚ�?             2@        ������������������������       �                     @        ^       a                   @H@���!pc�?             &@        _       `                 0c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        b       e                    �?؇���X�?             @        c       d                   �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        g       �                     �?��6}��?&            �N@       h       u                   �>@Ȩ�I��?#            �J@        i       t                 `fF<@և���X�?             5@       j       s                   �K@�q�q�?
             2@       k       r                   @G@���Q��?             $@       l       m                 03k:@և���X�?             @        ������������������������       �                     �?        n       o                 �|�<@�q�q�?             @        ������������������������       �                     �?        p       q                 X��B@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        v       �                    �?     ��?             @@       w       z                 ��9L@�>4և��?             <@       x       y                   �;@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        {       |                 `f�N@X�<ݚ�?             "@        ������������������������       �                      @        }       �                   �G@����X�?             @       ~       �                   �D@r�q��?             @              �                 X��@@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �@@      �?              @        ������������������������       �                     @        �       �                   �>@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�"�
�?�            0x@        �       �                    �?�D}1o��?K             `@       �       �                 �̌@�X����?5             V@        �       �                 P�@6YE�t�?            �@@        �       �                    �?�q�q�?             "@        ������������������������       �                     @        �       �                 �|Y:@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                 �|Y;@�8��8��?             8@       �       �                   �7@8�Z$���?	             *@       �       �                    �?�8��8��?             (@        ������������������������       �                      @        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 @33"@<|ۤ$�?             �K@        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?             H@        �       �                    �?z�G�z�?	             4@       �       �                    �?�	j*D�?             *@        �       �                   �-@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    &@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @      �?             <@        ������������������������       �                      @        �       �                 ���1@��
ц��?             :@       �       �                   �"@ҳ�wY;�?
             1@        ������������������������       �                     @        �       �                    �?և���X�?	             ,@       �       �                  �m#@�q�q�?             (@        ������������������������       �                     �?        �       �                 �[$@���!pc�?             &@        ������������������������       �                      @        �       �                 ��&@�q�q�?             "@        ������������������������       �                     �?        �       �                 @3�/@      �?              @        ������������������������       �                     @        �       �                   �0@���Q��?             @       �       �                 �|�;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �>@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                 �̼6@���?            �D@        �       �                   �/@�q�q�?             "@        �       �                 �|Y7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @      �?             @@       �       �                    @ �q�q�?             8@        �       �                 ��T?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        �       �                    �?      �?              @        ������������������������       �                      @        �       �                   @C@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �?�@��ED���?�             p@       �       �                   �8@X�GP>��?W            �_@        �       �                    �?$G$n��?            �B@        �       �                 ���@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���@�g�y��?             ?@        �       �                 ���@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     8@        �       �                    �?����?�?>            �V@        �       �                  ��@�7��?            �C@       ������������������������       �                     5@        �       �                 P�J@�����H�?             2@       �       �                 X�I@�C��2(�?             &@       ������������������������       �      �?              @        ������������������������       �                     @        �       �                 �|Y=@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        "            �I@        �       �                   �4@p6��%�?V            ``@        �       �                 03�0@f�Sc��?"            �H@       �       �                    �?և���X�?             <@        ������������������������       �                     @        �       �                    �?      �?             8@       �       �                 0S5 @���Q��?             4@        �       �                 @3�@���!pc�?             &@        ������������������������       ����Q��?             @        �       �                   �3@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             "@        ������������������������       �                     @        �       �                    �?�����?             5@       ������������������������       �        	             ,@        �       �                    @����X�?             @        �       �                     @      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �                       @3�@����!�?4            �T@        �       �                    :@�n_Y�K�?             *@        ������������������������       �                      @                                 �?@�eP*L��?             &@        ������������������������       �                      @                                �A@�q�q�?             "@        ������������������������       �z�G�z�?             @        ������������������������       �      �?             @              (                   �?�~t��?-            @Q@                             ��) @��hJ,�?,             Q@        ������������������������       �                     9@                                 �?>��C��?            �E@        	                      �|Y?@r�q��?
             (@       
                         �?�<ݚ�?             "@                              �|Y<@      �?             @        ������������������������       �                      @                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                `3@z�G�z�?             @        ������������������������       �                     @                              03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                              pf� @r֛w���?             ?@        ������������������������       �                     @              '                   �?�>4և��?             <@             &                  �?@���B���?             :@             %                �|�=@     ��?             0@                             @3�!@������?
             .@                              �|Y<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �<@r�q��?             (@        ������������������������       �                     @        !      "                ���"@�q�q�?             @        ������������������������       �                      @        #      $                �|Y=@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0M)KK��h2h3h4hVh<�h=Kub������������|d�_Z�?�7s@K�?��8��8�?9��8���?�&!��ȩ?��]tc�?F]t�E�?]t�E�?      �?      �?���Q��?)\���(�?�؉�؉�?ى�؉��?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�A�A�?��-��-�?              �?F]t�E�?�.�袋�?              �?�������?ffffff�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ����?����Ǐ�?              �?�?�������?              �?�������?�������?      �?                      �?���	A�?��	A���?UUUUUU�?UUUUUU�?A��)A�?�־a�?      �?        x6�;��?AL� &W�?qG�w��?w�qGܱ?      �?        n۶m۶�?�$I�$I�?�������?333333�?      �?      �?n۶m۶�?�$I�$I�?              �?      �?              �?        UUUUUU�?UUUUUU�?��y��y�?�a�a�?      �?        �q�q�?�q�q�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        a����?�{a���?      �?        ۶m۶m�?�$I�$I�?              �?      �?        �N̓��?��be�F�?��(\���?{�G�z�?�-��-��?�A�A�?�m۶m��?�$I�$I�?�$I�$I�?۶m۶m�?;�;��?ى�؉��?              �?UUUUUU�?UUUUUU�?              �?�������?�������?9��8���?�q�q�?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?      �?              �?      �?              �?              �?              �?      �?              �?      �?              �?                      �?      �?        �q�q�?r�q��?              �?F]t�E�?t�E]t�?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        �!XG��?;ڼOq��?+�R��?�	�[���?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?�������?333333�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?�$I�$I�?�m۶m��?�5��P�?(�����?              �?      �?        r�q��?�q�q�?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?              �?      �?      �?        333333�?�������?              �?      �?              �?        ���H���?�dxn�0�?QW�uE�?W�uE]�?]t�E]�?�E]t��?e�M6�d�?'�l��&�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?��7�}��?��)A��?�m۶m��?�$I�$I�?              �?      �?              �?      �?�������?�������?;�;��?vb'vb'�?333333�?�������?      �?                      �?      �?      �?              �?      �?                      �?      �?      �?              �?�;�;�?�؉�؉�?�������?�������?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        t�E]t�?F]t�E�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?�������?333333�?      �?      �?      �?                      �?              �?      �?        �q�q�?�q�q�?      �?                      �?28��1�?8��18�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?              �?      �?              �?      �?        �'�	�?��=aO��?����x<�?���p8�?к����?���L�?UUUUUU�?UUUUUU�?              �?      �?        ��{���?�B!��?۶m۶m�?�$I�$I�?      �?                      �?      �?        ��I��I�?l�l��?��[��[�?�A�A�?      �?        �q�q�?�q�q�?]t�E�?F]t�E�?      �?      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?        ��0�]��?BJ�eD�?����>�?������?۶m۶m�?�$I�$I�?              �?      �?      �?333333�?�������?t�E]t�?F]t�E�?�������?333333�?UUUUUU�?�������?              �?      �?              �?                      �?=��<���?�a�a�?      �?        �m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        %jW�v%�?jW�v%j�?;�;��?ى�؉��?      �?        t�E]t�?]t�E�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?�s��\�?)�3J���?KKKKKK�?�������?      �?        $�;��?qG�w��?�������?UUUUUU�?9��8���?�q�q�?      �?      �?      �?              �?      �?      �?                      �?�������?�������?      �?              �?      �?              �?      �?              �?        ���{��?�B!��?              �?�$I�$I�?�m۶m��?��؉���?ى�؉��?      �?      �?wwwwww�?�?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�)�rhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       T                    �?"��p�?�           8�@                                    @l��=���?�            p@                                  :@���۟�?P            `a@                                   �?��d��?            �O@        ������������������������       �                     $@                                    �?r�����?            �J@        ������������������������       �                      @                                   L@��x_F-�?            �I@       	                          �;@ZՏ�m|�?            �H@        
                           �?�q�q�?
             5@                                 �6@j���� �?             1@       ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     @                                  �8@h�����?             <@       ������������������������       �                     8@                                  �E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        1             S@               %                    �?vs�G��?L            �]@                                   �?�㙢�c�?             G@                                  �?�FVQ&�?            �@@                                ���,@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ;@                                �*%@��
ц��?             *@        ������������������������       �                     @               $                  18@�z�G��?             $@               #                 83�0@�<ݚ�?             "@        !       "                   �8@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        &       I                   @1@      �?3             R@       '       (                   �1@v ��?             �E@        ������������������������       �                     @        )       H                    �?X�<ݚ�?             B@       *       E                    �?j���� �?             A@       +       D                 ��Y.@���Q��?             >@       ,       -                   �5@�q�q�?             ;@        ������������������������       �                     @        .       9                   �@և���X�?             5@        /       8                 �&B@�q�q�?             "@       0       5                 ���@և���X�?             @        1       2                 ���@      �?             @        ������������������������       �                     �?        3       4                 �|Y:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        6       7                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        :       A                 ��&@      �?
             (@       ;       <                   �9@z�G�z�?             $@        ������������������������       �                     @        =       >                 �?�@�q�q�?             @        ������������������������       �                      @        ?       @                 @3�@      �?             @        ������������������������       �                      @        ������������������������       �                      @        B       C                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        F       G                   �;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        J       K                    �?\-��p�?             =@        ������������������������       �                     @        L       O                    @�㙢�c�?             7@        M       N                 ��T?@      �?             @       ������������������������       �                     @        ������������������������       �                     @        P       S                    �?�IєX�?             1@        Q       R                 �|Y>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             ,@        U       �                 ��D:@ҔOl�?!           `|@       V       [                    ,@t���|�?�            �t@        W       Z                    �?�8��8��?             (@        X       Y                    '@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        \       ]                     �?,_ʯ08�?�            �s@        ������������������������       �                      @        ^       o                    �?(�����?�            `s@        _       l                    �?�MI8d�?            �B@       `       a                     @�t����?             A@        ������������������������       �                     @        b       k                 �0@�r����?             >@       c       j                 �|Y=@@4և���?             <@        d       i                    <@�q�q�?             @       e       f                 �{@z�G�z�?             @        ������������������������       �                      @        g       h                 H�%@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                      @        m       n                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        p       �                   @@@($�pa�?�            q@       q       �                    �?�M��?|            �i@       r       �                   �+@�j�zZ��?y             i@       s       ~                     @lO�o���?k            �e@        t       u                    @V�a�� �?             =@        ������������������������       �                     @        v       y                   �'@�+e�X�?             9@        w       x                    5@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        z       {                 �|Y<@      �?             0@       ������������������������       �                     "@        |       }                 �|�=@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @               �                 �Y�@������?X             b@        �       �                    �?��?^�k�?            �A@        ������������������������       �                      @        �       �                    7@ 7���B�?             ;@        ������������������������       �                     *@        �       �                   �8@@4և���?             ,@        �       �                 `fF@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?lGts��?G            �[@        �       �                 ��(@r�q��?             (@       �       �                 �|Y=@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        �       �                 �|�=@ i���t�??            �X@       �       �                 �|Y=@`��F:u�?9            �U@       �       �                   �0@ ������?(            �O@        �       �                 pf�@z�G�z�?             @        ������������������������       �                     @        �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        %             M@        �       �                 ��) @      �?             8@       �       �                  sW@���N8�?             5@        ������������������������       ��q�q�?             @        ������������������������       �                     2@        �       �                 �̜!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �?�@�eP*L��?             &@        �       �                   �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��l!@z�G�z�?             @       �       �                   �?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ;@        ������������������������       �                     @        �       �                   �D@ ��ʻ��?/             Q@       ������������������������       �                     E@        �       �                 `f�)@ ��WV�?             :@       ������������������������       �                     2@        �       �                   �*@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03#?@Z��Yo��?O             _@        �       �                    �?�q�q�?             B@       �       �                  I>@     ��?             @@       �       �                     �?
j*D>�?             :@       �       �                   �J@���Q��?             9@       �       �                 03k:@�z�G��?             4@        ������������������������       �                     @        �       �                 ��=@ҳ�wY;�?
             1@       �       �                 �|�?@      �?             $@        ������������������������       �                     @        �       �                   `G@r�q��?             @       �       �                 `f�;@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y=@؇���X�?             @        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �Q@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 0�"K@N�zv�?9             V@        �       �                    @���H��?             E@        �       �                     @և���X�?             @        ������������������������       �                      @        �       �                 ���A@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                     �?��?^�k�?            �A@       �       �                 �|�<@ �q�q�?             8@        �       �                 `f�D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             4@        ������������������������       �                     &@        �       �                 03c@\X��t�?              G@       �       �                    �?      �?             B@        �       �                    �?p�ݯ��?             3@       �       �                   �8@      �?             (@        ������������������������       �                      @        �       �                   �H@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                 ��UO@և���X�?             @        ������������������������       �                      @        �       �                    �?���Q��?             @        �       �                    B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��#[@ҳ�wY;�?             1@       �       �                 �TL@������?             .@        ������������������������       �                     @        �       �                    �?�q�q�?             (@       �       �                     @�z�G��?	             $@       �       �                 `f�N@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ;@���Q��?             @        ������������������������       �                     �?        �       �                 �|�>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��R@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 @�:x@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������J54v��?l�����?�`�`�`�?�'�'�'�?����j�?��a����?EQEQ�?��뺮��?              �?�V�9�&�?Dj��V��?              �?�?�������?9/����?�>4և��?UUUUUU�?UUUUUU�?ZZZZZZ�?�������?              �?      �?                      �?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?              �?                      �?�N��?���؊��?d!Y�B�?�7��Mo�?|���?>����?UUUUUU�?UUUUUU�?              �?      �?                      �?�؉�؉�?�;�;�?      �?        333333�?ffffff�?�q�q�?9��8���?      �?      �?              �?      �?                      �?      �?              �?      �?qG�w��?G�w��?              �?r�q��?�q�q�?�������?ZZZZZZ�?333333�?�������?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?              �?      �?                      �?      �?      �?              �?      �?                      �?a����?�{a���?      �?        �7��Mo�?d!Y�B�?      �?      �?      �?                      �?�?�?UUUUUU�?UUUUUU�?      �?                      �?      �?        z\��W&�?�$�f�?j�ƀi�?��?����?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?����6b�?��J�?      �?        Q���P�?y�W�x�?��L���?L�Ϻ��?<<<<<<�?�?      �?        �������?�?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?~ڧ}ڧ�?,�,��?	݋н�?��{��?/�Q����?��s��2�?�Ȥx��?�C��:��?��{a�?a���{�?      �?        R���Q�?���Q��?9��8���?�q�q�?              �?      �?              �?      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?        ��y�!�?C:o1��?_�_��?�A�A�?      �?        	�%����?h/�����?      �?        n۶m۶�?�$I�$I�?      �?      �?              �?      �?              �?        �<%�S��?�־a�?�������?UUUUUU�?/�袋.�?F]t�E�?              �?      �?              �?        /�����?����X�?�u�7[��?Ȥx�L��?��}��}�?AA�?�������?�������?      �?              �?      �?              �?      �?              �?              �?      �?��y��y�?�a�a�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ]t�E�?t�E]t�?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        �������?�?      �?        O��N���?;�;��?      �?              �?      �?              �?      �?        !�B!�?���{��?�������?�������?      �?      �?;�;��?b'vb'v�?�������?333333�?333333�?ffffff�?              �?�������?�������?      �?      �?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?�������?�������?      �?                      �?      �?                      �?      �?        颋.���?/�袋.�?�0�0�?��y��y�?۶m۶m�?�$I�$I�?              �?333333�?�������?              �?      �?        _�_��?�A�A�?�������?UUUUUU�?      �?      �?              �?      �?              �?              �?        !Y�B�?��Moz��?      �?      �?Cy�5��?^Cy�5�?      �?      �?      �?        �������?�������?              �?      �?        �$I�$I�?۶m۶m�?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �������?�������?wwwwww�?�?      �?        UUUUUU�?UUUUUU�?ffffff�?333333�?�������?�������?              �?      �?        333333�?�������?              �?      �?      �?      �?                      �?      �?      �?      �?                      �?              �?�������?�������?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJX"4qhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       L                    �?|��;;��?�           8�@                                   �?g�R��?y            �g@                                   &@�C��2(�?1            @S@                                ���,@      �?             @        ������������������������       �                     �?                                `�@1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        	                           �?���;QU�?.            @R@       
                            �?P����?'            �M@                                   �?�nkK�?             7@                               ��A@���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                      @        ������������������������       �                     B@                                �|Y=@����X�?             ,@        ������������������������       �                     @                                     @      �?              @        ������������������������       �                     @                                 S�2@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                ���@
�ۓQ{�?H            @\@                                03S@��S�ۿ?             .@        ������������������������       �                      @                                �|�9@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@               A                    �?~���L0�?@            �X@              .                 �|Y=@���+�?1            �R@                +                  �}S@��Q��?             4@       !       *                    �?      �?	             0@       "       #                      @������?             .@        ������������������������       �                     @        $       %                    7@���Q��?             $@        ������������������������       �                     @        &       )                 �0@�q�q�?             @       '       (                   �<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ,       -                   �8@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        /       8                    C@PN��T'�?%             K@       0       7                 ��(@@4և���?             E@        1       6                 �|�=@r�q��?             2@       2       3                    �?@�0�!��?             1@        ������������������������       ��q�q�?             @        4       5                 ���@؇���X�?	             ,@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     8@        9       :                  �>@�q�q�?             (@        ������������������������       �                     @        ;       @                    N@      �?              @       <       ?                   @G@����X�?             @       =       >                   @N@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        B       C                 �n6@      �?             8@        ������������������������       �                     @        D       K                 @��v@���y4F�?             3@       E       F                    �?r�q��?             2@        ������������������������       �                      @        G       J                    6@      �?
             0@        H       I                  D�Q@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        M       �                    �?`� w���?F           H�@        N       k                     @ ��3j�?o             f@       O       Z                   �B@�:�H:�?@            @[@       P       Y                    �?��pBI�?-            @R@       Q       X                   �7@�7��?            �C@        R       W                   �;@�t����?             1@        S       T                   �6@����X�?             @        ������������������������       �                     @        U       V                   �'@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     6@        ������������������������       �                     A@        [       j                    �?      �?             B@       \       c                   �*@      �?             8@        ]       ^                    D@��
ц��?             *@        ������������������������       �                     @        _       b                   �'@      �?              @       `       a                   �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        d       e                     �?"pc�
�?             &@        ������������������������       �                     @        f       g                   �E@�q�q�?             @        ������������������������       �                     @        h       i                   @F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        l       �                    �?ҳ�wY;�?/             Q@       m       p                    @      �?              E@        n       o                 @3�2@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        q       �                    �?X�<ݚ�?             B@       r                          �9@��
ц��?             :@       s       z                   �3@�n_Y�K�?             *@        t       y                 `F�+@�q�q�?             @       u       x                 �&B@z�G�z�?             @        v       w                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        {       |                   �6@؇���X�?             @        ������������������������       �                     @        }       ~                 @3�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03�1@�	j*D�?
             *@       �       �                   �D@"pc�
�?	             &@       �       �                 P��@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �>@z�G�z�?             $@       �       �                   �;@�����H�?             "@        �       �                   �1@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                  `/@ȵHPS!�?             :@        ������������������������       �                     �?        �       �                 ��T?@HP�s��?             9@       ������������������������       �                     1@        �       �                 ��p@@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                    #@�b��R��?�            �u@        �       �                     @�q�q�?             8@        ������������������������       �                     &@        �       �                    @��
ц��?
             *@        �       �                    �?r�q��?             @       �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @����X�?             @        ������������������������       �                     �?        �       �                 `f�9@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 `ff:@(\�����?�             t@       �       �                   @E@�m(�X�?�            �o@       �       �                 �?�@�q����?�            �k@        �       �                     @ qP��B�?9            �U@        ������������������������       �        	             *@        �       �                   �7@��pBI�?0            @R@        ������������������������       �                     7@        �       �                   �8@`2U0*��?"             I@        �       �                 `fF@z�G�z�?             @        �       �                 �&b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y=@����?�?            �F@        ������������������������       �                     3@        �       �                 �|Y>@ ��WV�?             :@       �       �                  sW@��S�ۿ?             .@       �       �                 pf�@      �?              @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     &@        �       �                 �|�=@����&�?T            �`@       �       �                    &@����"$�?:            �U@       �       �                 ��) @X�;�^o�?%            �K@        �       �                   �4@�����H�?             ;@        �       �                   �3@�q�q�?             "@       �       �                   �1@���Q��?             @        ������������������������       ��q�q�?             @        ������������������������       �      �?              @        �       �                 @3�@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �        
             2@        �       �                   �<@؇���X�?             <@       �       �                     @���}<S�?             7@        �       �                    5@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                 @�!@      �?
             0@        �       �                   �:@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y=@���Q��?             @       �       �                 ���"@�q�q�?             @        ������������������������       �                     �?        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ?@        �       �                     @      �?             H@        �       �                   �3@�<ݚ�?
             2@       �       �                    @@���|���?             &@        ������������������������       �                     @        �       �                   @B@�q�q�?             @        ������������������������       �                     @        �       �                   @D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ?@������?             >@        �       �                 �̌!@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 pf� @���B���?             :@        �       �                   �A@X�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �����X�?             @        ������������������������       �        
             1@        ������������������������       �                    �A@        �       �                   �>@�	j*D�?%            @P@        �       �                    �?�q�q�?             5@       �       �                 X��A@�d�����?             3@        ������������������������       �                     @        �       �                     �?�n_Y�K�?             *@       �       �                   �F@�q�q�?             (@        ������������������������       �                      @        �       �                   `G@���Q��?             $@        ������������������������       �                      @        �       �                 `fF<@      �?              @       �       �                    M@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       
                    @��2(&�?             F@       �                       ��#[@ >�֕�?            �A@       �                          �?      �?             @@                                �C@�g�y��?             ?@       ������������������������       �                     1@                                �E@@4և���?             ,@                               x#J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?              	                X��C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?X�<ݚ�?             "@                              �|�;@z�G�z�?             @        ������������������������       �                     @                              �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������|d�_Z�?�7s@K�?��sK���?+Fڱ�?F]t�E�?]t�E�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�1bĈ�?�ܹs���?'u_[�?�V'u�?d!Y�B�?�Mozӛ�?�a�a�?��y��y�?      �?                      �?              �?              �?�$I�$I�?�m۶m��?              �?      �?      �?              �?�������?�������?      �?                      �?2�s�8�?��Ź��?�������?�?      �?        �؉�؉�?;�;��?              �?      �?        ����>4�?������?�n0E>��?�"�u�)�?ffffff�?�������?      �?      �?�?wwwwww�?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?              �?      �?      �?      �?                      �?&���^B�?h/�����?n۶m۶�?�$I�$I�?�������?UUUUUU�?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?              �?        �������?�������?      �?              �?      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?              �?      �?              �?6��P^C�?(������?�������?UUUUUU�?              �?      �?      �?�������?�������?      �?                      �?      �?                      �?�|r���?c��?j�`���?K�O�v�?\����չ?Ṷ�H��?����?���Ǐ�?�A�A�?��[��[�?�?<<<<<<�?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?                      �?              �?              �?      �?      �?      �?      �?�;�;�?�؉�؉�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?      �?UUUUUU�?�������?              �?      �?        r�q��?�q�q�?�؉�؉�?�;�;�?;�;��?ى�؉��?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        ;�;��?vb'vb'�?F]t�E�?/�袋.�?�������?�������?      �?                      �?      �?              �?        �������?�������?�q�q�?�q�q�?      �?      �?      �?                      �?      �?                      �?��N��N�?�؉�؉�?              �?q=
ףp�?{�G�z�?      �?              �?      �?              �?      �?        ��)kʚ�?eMYS֔�?�������?�������?              �?�;�;�?�؉�؉�?�������?UUUUUU�?      �?      �?      �?                      �?      �?        �$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?        fffff��?ffffff�?]]]]]]�?�?� O	��?pX���o�?��}A�?�}A_З?      �?        ���Ǐ�?����?      �?        ���Q��?{�G�z�?�������?�������?      �?      �?      �?                      �?      �?        ��I��I�?l�l��?      �?        O��N���?;�;��?�������?�?      �?      �?      �?              �?      �?      �?              �?        �Dz�rv�?��~5&�?YS֔5e�?6eMYSִ?�־a��?J��yJ�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?        ۶m۶m�?�$I�$I�?ӛ���7�?d!Y�B�?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?�������?�������?      �?                      �?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?      �?              �?      �?              �?              �?      �?9��8���?�q�q�?]t�E]�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        wwwwww�?�?      �?      �?      �?                      �?��؉���?ى�؉��?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?      �?              �?        vb'vb'�?;�;��?UUUUUU�?UUUUUU�?y�5���?Cy�5��?              �?ى�؉��?;�;��?UUUUUU�?UUUUUU�?              �?�������?333333�?      �?              �?      �?�������?333333�?              �?      �?                      �?      �?              �?        ��.���?t�E]t�?��+��+�?�A�A�?      �?      �?��{���?�B!��?      �?        n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?r�q��?�q�q�?�������?�������?              �?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ;�3whG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       l                    �?�����?�           8�@               M                    �?�^� ���?�            �m@              L                 03[=@�Q@�d�?�            �g@              K                 03�;@栤k��?W             _@              B                 Ь�9@��[�A�?V            �^@              1                    �?xZ�l ��?J            �Z@                                  �?Gq����?9            @U@                                  �-@ 	��p�?             =@        	       
                 H�%@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     :@               ,                 03�0@��>4և�?(             L@              #                 �|�=@�J��%�?#            �H@                               `fV$@�P�*�?             ?@                               @3�@ҳ�wY;�?             1@                                 �3@�q�q�?             "@        ������������������������       �                     �?                                P�@      �?              @                               �|�;@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                  �9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                 ��-@؇���X�?	             ,@                               `f�)@�8��8��?             (@       ������������������������       �                     @                                   :@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        !       "                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        $       )                     @r�q��?             2@       %       (                   �'@�C��2(�?	             &@        &       '                   �J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        *       +                   �C@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        -       0                     @؇���X�?             @        .       /                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        2       3                 P��%@���|���?             6@        ������������������������       �                      @        4       5                     @�z�G��?             4@        ������������������������       �                     @        6       9                    �?      �?             0@        7       8                    @      �?              @        ������������������������       �                     @        ������������������������       �                     @        :       ;                    @      �?              @        ������������������������       �                     @        <       =                    @���Q��?             @        ������������������������       �                     �?        >       ?                 �|Y<@      �?             @        ������������������������       �                      @        @       A                  ��6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        C       D                     �?��S�ۿ?             .@        ������������������������       �                     �?        E       J                    :@@4և���?             ,@       F       I                    �?ףp=
�?             $@       G       H                   �E@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        *             P@        N       c                 �|�:@ڡR����?            �H@       O       X                 03�;@      �?             @@        P       Q                     @�����H�?	             2@       ������������������������       �                     $@        R       S                    @      �?              @        ������������������������       �                     @        T       W                    @���Q��?             @       U       V                 ��l4@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        Y       `                    1@և���X�?
             ,@       Z       [                 ��T?@      �?              @        ������������������������       �                     @        \       ]                    �?      �?             @        ������������������������       �                     �?        ^       _                    %@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        a       b                      @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        d       e                     @�t����?             1@        ������������������������       �                     @        f       g                    @$�q-�?             *@       ������������������������       �                     $@        h       k                    @�q�q�?             @       i       j                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        m       �                     �?h��Z }�?$           �}@        n       s                   �:@Bԅ���?7            �W@        o       p                 �U�X@�C��2(�?             &@       ������������������������       �                      @        q       r                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        t       �                   �J@0,Tg��?2             U@       u       �                   `A@d��0u��?$             N@       v       �                    @@��S���?             >@       w       x                    �?      �?
             0@        ������������������������       �                     @        y       z                    <@�	j*D�?             *@        ������������������������       �                     �?        {       |                 �|Y=@      �?             (@        ������������������������       �                      @        }       ~                 `fF<@�z�G��?             $@        ������������������������       �                     @               �                   �>@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?؇���X�?	             ,@        ������������������������       �                      @        �       �                 ��I*@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        �       �                   �G@z�G�z�?             >@       �       �                 �|Y<@�LQ�1	�?             7@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?ףp=
�?
             4@        ������������������������       �                     @        �       �                 �|Y>@؇���X�?             ,@        ������������������������       �                      @        �       �                 0��J@�q�q�?             @        ������������������������       �                     @        �       �                   @A@�q�q�?             @        ������������������������       �                     �?        �       �                 ��n^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �H@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     8@        �       �                    �?�%F@ ��?�            �w@       �       �                     @������?�             t@        �       �                   �*@@݈g>h�?.             S@       �       �                    @�:pΈ��?             I@        ������������������������       �                     @        �       �                 ��Y)@��0{9�?            �G@        �       �                    5@�t����?             1@        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        ������������������������       �                     &@        �       �                 �|�<@r�q��?             >@        ������������������������       �                     ,@        �       �                 �|�=@     ��?	             0@        ������������������������       �                     �?        �       �                    @@������?             .@        ������������������������       �                     @        �       �                   �A@�q�q�?             (@        ������������������������       �                      @        �       �                   @D@z�G�z�?             $@        ������������������������       �                     @        �       �                    G@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     :@        �       �                 �T)D@��w��?�            �n@       �       �                    �?�l�T{�?�             n@        �       �                    7@��S�ۿ?             >@        ������������������������       �                      @        ������������������������       �                     <@        �       �                   @@@�S	���?�            `j@       �       �                 ���#@ �Cc}�?j             e@       �       �                    �?H%u��?_            �b@        �       �                 �|Y=@�LQ�1	�?             7@        �       �                    ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                  s�@ףp=
�?             4@        ������������������������       �                     @        �       �                 ��(@؇���X�?	             ,@       ������������������������       �8�Z$���?             *@        ������������������������       �                     �?        �       �                 �|�=@X�GP>��?P            �_@       �       �                   �<@8@W"�h�?M            @^@       �       �                 �?�@ ,U,?��?4            �T@       �       �                 ���@���J��?            �I@        �       �                 ���@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                    �D@        �       �                 0S5 @      �?             @@        �       �                 @3�@      �?	             (@        �       �                   �4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        �       �                   �5@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                   �:@P���Q�?             4@       ������������������������       �        
             0@        �       �                   �;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y=@�?�'�@�?             C@        �       �                 ���"@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                  sW@(N:!���?            �A@        �       �                 pf�@�q�q�?             "@       ������������������������       �                     @        ������������������������       ����Q��?             @        �       �                 ��) @ ��WV�?             :@       ������������������������       �                     7@        �       �                 pf� @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 P�@r�q��?             @        ������������������������       �                     @        �       �                    ?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                    �E@        �       �                    ;@���Q��?             @        ������������������������       �                      @        �       �                 �|�>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �                            @p�ݯ��?%            �L@        �       �                    �?      �?	             0@        �       �                    *@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    :@X�Cc�?             ,@       �       �                    �?"pc�
�?             &@       �       �                   @.@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @                                 #@���� �?            �D@                                �?\X��t�?             7@        ������������������������       �                      @                                 �?�ՙ/�?             5@        ������������������������       �                     @                              ���A@և���X�?
             ,@                             @3�4@�����H�?             "@       ������������������������       �                     @        	      
                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?�X�<ݺ?             2@                              �|Y7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�����������������?��܍��?��"`c��?�[�'��?�٨�l��?����
�?B!��?��{���?�:ڼO�?z��!X�?�+J�#�?�w�Zn�?�?�������?�{a���?������?UUUUUU�?UUUUUU�?              �?      �?                      �?I�$I�$�?۶m۶m�?9/����?c}h���?�Zk����?�RJ)���?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?�������?              �?      �?              �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?      �?      �?                      �?UUUUUU�?�������?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?�m۶m��?              �?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        F]t�E�?]t�E]�?      �?        333333�?ffffff�?              �?      �?      �?      �?      �?              �?      �?              �?      �?              �?�������?333333�?      �?              �?      �?              �?      �?      �?              �?      �?        �?�������?              �?�$I�$I�?n۶m۶�?�������?�������?�q�q�?�q�q�?              �?      �?                      �?              �?      �?                      �?����X�?����S��?      �?      �?�q�q�?�q�q�?              �?      �?      �?              �?�������?333333�?      �?      �?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?      �?        �������?�������?              �?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        vr.�e�?)6F�i�?�S��8�?�X�0Ҏ�?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?                      �?�y��y��?1�0��?DDDDDD�?wwwwww�?�������?�?      �?      �?      �?        vb'vb'�?;�;��?              �?      �?      �?      �?        ffffff�?333333�?      �?        �������?333333�?              �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?�������?      �?                      �?�������?�������?��Moz��?Y�B��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?        :��|���?�(j9�?c��*��?�싨�ٷ?�P^Cy�?Cy�5��?��Q���?�Q����?      �?        m�w6�;�?L� &W�?<<<<<<�?�?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?        �������?UUUUUU�?      �?              �?      �?              �?wwwwww�?�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?        333333�?�������?      �?      �?      �?              �?        M!��?��~Y�?}*X}*X�?�>�>�?�������?�?              �?      �?        �ƴ	(E�?1�Y��ֵ?%I�$I��?۶m۶m�?)\���(�?���Q��?��Moz��?Y�B��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?        ۶m۶m�?�$I�$I�?;�;��?;�;��?      �?        ���p8�?����x<�?��#��Z�?�C��2(�?��ˊ��?��FS�׮?______�?�?�������?�������?      �?                      �?      �?              �?      �?      �?      �?�������?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?        ffffff�?�������?      �?              �?      �?              �?      �?        ������?y�5���?UUUUUU�?UUUUUU�?      �?                      �?|�W|�W�?�A�A�?UUUUUU�?UUUUUU�?      �?        �������?333333�?O��N���?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?^Cy�5�?Cy�5��?      �?      �?      �?      �?              �?      �?        �m۶m��?%I�$I��?F]t�E�?/�袋.�?�������?�������?      �?                      �?      �?              �?        jW�v%j�?,Q��+�?!Y�B�?��Moz��?              �?�<��<��?�a�a�?      �?        ۶m۶m�?�$I�$I�?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��8��8�?�q�q�?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�3hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       d                    �?�E	�rQ�?�           8�@               Y                   XB@@�h�|5�?�            �p@              R                 03#?@>�V�n��?q             g@                                  @.��|\�?j            �e@        ������������������������       �                     ,@               ;                    �?��Y���?b            �c@                                    @�k��(A�?H            �]@                                  �H@ s�n_Y�?              J@       	                          �6@,���i�?            �D@       
                          `2@"pc�
�?             6@                                 �B@�X�<ݺ?             2@       ������������������������       �                     ,@                                  �C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   ?@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                 	<@�}�+r��?             3@                                  D@@4և���?	             ,@       ������������������������       �                     $@                                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                    �?�eP*L��?             &@                                ���;@      �?              @        ������������������������       �                     @        ������������������������       �                     @                                   L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        !       *                    �?҄��?(            �P@        "       %                 ���@4?,R��?             B@        #       $                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        &       '                 ���,@�C��2(�?            �@@       ������������������������       �                     6@        (       )                  S�-@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        +       ,                 ���@���Q��?             >@        ������������������������       �                     @        -       4                 �|Y>@ �o_��?             9@       .       /                   �5@z�G�z�?             4@        ������������������������       �                     @        0       1                  sW@      �?	             0@        ������������������������       �                      @        2       3                 ��*@؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @        5       :                 ��Y.@���Q��?             @       6       7                 ��n @�q�q�?             @        ������������������������       �                     �?        8       9                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        <       =                    '@H�z�G�?             D@        ������������������������       �                     @        >       A                   �;@      �?             A@        ?       @                    �?r�q��?	             (@        ������������������������       �                      @        ������������������������       �                     $@        B       K                    D@�X����?             6@       C       J                    @@�0�!��?
             1@       D       G                    �?z�G�z�?	             .@       E       F                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        H       I                 �|Y=@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        L       Q                   �H@z�G�z�?             @       M       N                   �E@�q�q�?             @        ������������������������       �                     �?        O       P                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        S       T                    �?�θ�?             *@        ������������������������       �                     �?        U       V                 ��T?@r�q��?             (@        ������������������������       �                     @        W       X                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        Z       c                 ���Q@0��P�?1            �T@        [       ^                 �|�:@�חF�P�?             ?@        \       ]                     @      �?	             0@       ������������������������       �                     .@        ������������������������       �                     �?        _       `                    �?������?
             .@       ������������������������       �                     "@        a       b                   �F@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �I@        e       r                    @�,���?           �{@        f       g                     @�z�G��?	             4@        ������������������������       �                     @        h       m                    �?ҳ�wY;�?             1@       i       l                    @X�<ݚ�?             "@       j       k                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        n       q                     @      �?              @       o       p                 pf�@@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        s       �                     �?x���L��?           �z@        t       �                   �J@2E�=<��?>            �X@       u       �                    �?H���I�?2            �S@        v       �                    �?��S���?             >@       w       �                  �}S@���Q��?             9@       x       y                 �ܵ<@"pc�
�?             &@        ������������������������       �                     �?        z       {                 �|Y<@ףp=
�?             $@        ������������������������       �                     @        |                         �>@z�G�z�?             @        }       ~                 ��2>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 t�is@և���X�?             ,@       �       �                   �8@���!pc�?             &@        ������������������������       �                     @        �       �                   �H@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �7@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �>@ \� ���?             �H@        �       �                   �9@��.k���?             1@        ������������������������       �                     @        �       �                 `fF<@ףp=
�?             $@       �       �                    D@z�G�z�?             @        ������������������������       �                      @        �       �                   @G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��yC@     ��?             @@        �       �                 �|�<@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���[@�>����?             ;@       �       �                 `�iJ@���7�?             6@        �       �                  x#J@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        �       �                 ���a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                  Y>@�}�+r��?             3@        �       �                    �?r�q��?             @        ������������������������       �                     �?        �       �                   �Q@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        �       �                  ��@�Iy4�%�?�            `t@        �       �                 ���@0�z��?�?-             O@       ������������������������       �                     B@        �       �                   @4@ ��WV�?             :@        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        �       �                    0@Pe6�p�?�            �p@       �       �                   �0@2%ޑ��?�            @j@        �       �                    )@      �?              @        ������������������������       �                      @        �       �                 �̌!@�q�q�?             @       ������������������������       �z�G�z�?             @        ������������������������       �                     �?        �       �                 `�X.@(r3.��?~            @i@       �       �                   �@     ��?x             h@        �       �                   �<@�'�`d�?            �@@        ������������������������       �        	             $@        �       �                   @@@8����?             7@       �       �                    �?b�2�tk�?             2@       �       �                 �|Y=@d}h���?	             ,@        ������������������������       �                     �?        �       �                 ��(@8�Z$���?             *@       ������������������������       �r�q��?             (@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�J��_��?`            �c@        �       �                 �� @��S�ۿ?             .@       �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                     @�5?,R�?Y             b@        �       �                   @D@dP-���?            �G@       �       �                    &@�X�<ݺ?             B@        �       �                    5@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                 �|�<@���N8�?             5@       ������������������������       �        
             ,@        �       �                 �|�=@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    G@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?�$��y��?;            @X@       �       �                 �|�=@��a�n`�?9            @W@       �       �                 @3�@�nkK�?)            @Q@        ������������������������       �                     :@        �       �                 @3�!@Du9iH��?            �E@       �       �                   �:@      �?             8@       �       �                   �3@      �?
             0@        �       �                 pf� @z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 ��) @      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             3@        �       �                   �?@      �?             8@        �       �                   �>@�q�q�?             @       �       �                 (Se!@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    D@�����H�?             2@       �       �                   @C@"pc�
�?	             &@       �       �                   @@@ףp=
�?             $@       �       �                 �?�@r�q��?             @        ������������������������       �                     �?        �       �                 ��I @z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?���Q��?             $@        ������������������������       �                     @        �       �                 X�lA@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �                        �T�I@ 7���B�?!             K@       ������������������������       �                     H@                                 �?�q�q�?             @                                ;@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������JP���?7j_Q��?�E(B�?v�{��^�?�r�4�-�?�F��*i�?MYS֔5�?YS֔5e�?              �?-n����?�Ȟ��t�?~ylE�p�?A�Iݗ��?;�;��?�;�;�?8��18�?�����?F]t�E�?/�袋.�?�q�q�?��8��8�?              �?      �?      �?      �?                      �?      �?      �?      �?                      �?(�����?�5��P�?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?                      �?t�E]t�?]t�E�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        N6�d�M�?�d�M6��?r�q��?�8��8��?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?]t�E�?              �?t�E]t�?F]t�E�?      �?                      �?333333�?�������?              �?
ףp=
�?�Q����?�������?�������?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?ffffff�?333333�?      �?              �?      �?UUUUUU�?�������?      �?                      �?�E]t��?]t�E]�?ZZZZZZ�?�������?�������?�������?۶m۶m�?�$I�$I�?              �?      �?              �?      �?              �?      �?              �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?ى�؉��?�؉�؉�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        8��18�?���|�?��RJ)��?�Zk����?      �?      �?              �?      �?        �?wwwwww�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�$jN�?el��W��?333333�?ffffff�?              �?�������?�������?r�q��?�q�q�?�������?UUUUUU�?              �?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?W�9�&�?�&oe��?��>4և�?����S��?Q�Ȟ���?^-n����?�������?�?�������?333333�?F]t�E�?/�袋.�?      �?        �������?�������?              �?�������?�������?      �?      �?              �?      �?                      �?�$I�$I�?۶m۶m�?F]t�E�?t�E]t�?      �?              �?      �?              �?      �?                      �?�������?�������?              �?      �?        
^N��)�?և���X�?�?�������?      �?        �������?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?              �?              �?      �?      �?�������?�������?              �?      �?        �Kh/��?h/�����?�.�袋�?F]t�E�?�q�q�?�q�q�?      �?                      �?      �?        �������?�������?              �?      �?        �5��P�?(�����?�������?UUUUUU�?      �?        �������?�������?      �?                      �?      �?        2���\w�?n�
�E�?|���{�?�B!��?      �?        O��N���?;�;��?      �?      �?      �?                      �?      �?        �|���?���>��?�������?�A�A�?      �?      �?              �?UUUUUU�?UUUUUU�?�������?�������?      �?        &����?�g����?     ��?      �?6�d�M6�?'�l��&�?      �?        d!Y�B�?8��Moz�?�8��8��?9��8���?I�$I�$�?۶m۶m�?              �?;�;��?;�;��?�������?UUUUUU�?      �?                      �?      �?        d�^�.�?�%w��?�������?�?      �?      �?              �?      �?              �?        �q�q�?�q�q�?�����F�?W�+�ɵ?��8��8�?�q�q�?�������?�?              �?      �?        ��y��y�?�a�a�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        /�袋.�?F]t�E�?              �?      �?        ����?W?���?�s�9��?�c�1Ƹ?�Mozӛ�?d!Y�B�?      �?        qG�w��?w�qGܱ?      �?      �?      �?      �?�������?�������?      �?      �?      �?              �?              �?      �?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?              �?�q�q�?�q�q�?/�袋.�?F]t�E�?�������?�������?�������?UUUUUU�?      �?        �������?�������?      �?      �?      �?              �?                      �?      �?              �?        �������?333333�?      �?        �$I�$I�?۶m۶m�?              �?      �?        	�%����?h/�����?      �?        UUUUUU�?UUUUUU�?333333�?�������?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ� �NhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       Z                    �?�t����?�           8�@               I                 �|�=@�桐-�?�            @p@              H                 �̌R@�g�Ф��?q             f@                                  �?���-|$�?b            @c@                                   �?д>��C�?$             M@                                   @��p\�?            �D@        ������������������������       �                     "@               	                 �{&@     ��?             @@       ������������������������       �                     2@        
                         S�-@d}h���?             ,@                                �|Y6@      �?             @                                 �-@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                `�@1@j���� �?             1@                                   �?�<ݚ�?             "@                                  �?      �?              @        ������������������������       �                     @                                �|Y=@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @               A                 �|Y=@�q�Q�?>             X@              ,                   �3@��.���?6            �U@               #                    �?      �?             B@              "                 ��	6@���y4F�?             3@                                   @      �?              @        ������������������������       �                     �?                !                 `fF.@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        $       +                 03�=@�t����?             1@       %       *                    +@$�q-�?             *@       &       '                     @r�q��?             @       ������������������������       �                     @        (       )                 `f7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        -       4                     @���Q��?             I@        .       /                     �?P���Q�?             4@        ������������������������       �                     �?        0       3                   �9@�}�+r��?
             3@        1       2                   �+@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        5       8                    �?d��0u��?             >@       6       7                   �@���Q��?             4@        ������������������������       �                      @        ������������������������       �        	             (@        9       @                 ���9@�z�G��?             $@       :       ;                   �&@և���X�?             @        ������������������������       �                      @        <       ?                    �?���Q��?             @       =       >                   �;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        B       G                    �?z�G�z�?             $@        C       D                     @      �?             @        ������������������������       �                     �?        E       F                 pf�'@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        J       K                 ��n @�}#���?2            �T@        ������������������������       �                     �?        L       M                   @C@��p\�?1            �T@        ������������������������       �                     F@        N       Y                    @�S����?             C@       O       X                   �G@�����H�?             B@        P       W                     @���y4F�?
             3@       Q       V                    :@      �?	             0@        R       S                   �3@r�q��?             @        ������������������������       �                     @        T       U                   �E@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                      @        [       �                  x#J@���{.��?,           0|@       \       �                    �?|D�]�|�?           �x@       ]       z                    �?�H�KY�?�            Pu@        ^       i                 �|Y=@���5��?$            �L@        _       `                     �?����X�?
             ,@        ������������������������       �                     �?        a       h                 ��Y&@�θ�?	             *@       b       g                   @@      �?              @       c       d                 ���@����X�?             @        ������������������������       �                      @        e       f                   �5@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        j       q                   `A@Du9iH��?            �E@       k       p                     �?(;L]n�?             >@        l       o                 ��2>@      �?              @        m       n                 �ܵ<@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     6@        r       y                   �A@8�Z$���?	             *@       s       x                  �>@      �?              @       t       w                     �?؇���X�?             @        u       v                    <@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        {       �                     �?�
0����?�            �q@        |       �                   �G@      �?             F@       }       �                   �<@��G���?            �B@        ~                        `f�D@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��<:@��hJ,�?             A@        ������������������������       �                     ,@        �       �                    C@      �?             4@       �       �                   �>@�n_Y�K�?	             *@       �       �                 �|Y=@����X�?             @        ������������������������       �                     �?        �       �                 `fF<@r�q��?             @        �       �                 �|�?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `fF:@և���X�?             @        ������������������������       �                     �?        �       �                   �J@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�8��8��?�             n@        �       �                   `3@@4և���?             <@       �       �                  ��@ ��WV�?             :@        ������������������������       �                     @        �       �                   @'@P���Q�?             4@       �       �                 X��A@�X�<ݺ?             2@       ������������������������       �@4և���?	             ,@        ������������������������       �                     @        ������������������������       �                      @        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �>@��-#���?�            �j@       �       �                 �?�@���C�:�?e            `b@        ������������������������       �        -            �N@        �       �                   �+@X�EQ]N�?8            �U@       �       �                 @3�@     ��?,             P@        ������������������������       �      �?              @        �       �                     @���-T��?*             O@        �       �                 �|Y=@�S����?             3@       ������������������������       �                     &@        �       �                 �|�=@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �3@(L���?            �E@        �       �                 ��Y @���Q��?             $@        �       �                   �2@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                 pf� @�FVQ&�?            �@@        ������������������������       �                     1@        �       �                   �:@      �?             0@       ������������������������       �                     $@        �       �                   �;@�q�q�?             @        ������������������������       �                     �?        �       �                   �<@z�G�z�?             @        ������������������������       �                     @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        �       �                     @�?�<��?.            @P@        �       �                    F@�r����?             >@       �       �                 `fF)@"pc�
�?             6@        ������������������������       �                     @        �       �                   @A@������?	             1@        �       �                    1@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @D@8�Z$���?             *@       ������������������������       �                     "@        ������������������������       �      �?             @        ������������������������       �                      @        �       �                 @3�@(N:!���?            �A@       �       �                 �&B@�<ݚ�?             2@       ������������������������       �        	             (@        �       �                   �@�q�q�?             @        ������������������������       �                     �?        �       �                 �?�@���Q��?             @        ������������������������       �                     �?        �       �                   �?@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     1@        �       �                    @��U/��?&            �L@        �       �                     @      �?	             (@        ������������������������       �                     @        �       �                    �?և���X�?             @        �       �                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 pf�C@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     @:	��ʵ�?            �F@        ������������������������       �                     (@        �       �                    0@r٣����?            �@@        �       �                 �=/@���Q��?             $@       �       �                    �?և���X�?             @        ������������������������       �                      @        �       �                 P��)@z�G�z�?             @        �       �                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?���}<S�?             7@        ������������������������       �                     @        �       �                    '@ףp=
�?             4@        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    @      �?             @        ������������������������       �                     �?        �       �                 83�@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     .@        �       �                   �1@�F�j��?!            �J@        ������������������������       �                     @        �                           �?�[�IJ�?            �G@       �                         @I@��.k���?             A@       �                          �?��S���?             >@       �       �                  �}S@      �?             4@        ������������������������       �                     @        �                          ?@�θ�?	             *@       �                        �U�X@      �?              @        �       �                 0�HU@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                              �UcV@���Q��?             @        ������������������������       �                     �?                              @�ys@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                              �|Y>@���Q��?             $@        ������������������������       �                      @        	                      ���R@      �?              @       
                      03�M@�q�q�?             @                                G@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                              p�O@�	j*D�?             *@                             �|�>@      �?              @                                ;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������G�+J>�?r%�k���?[��Z���?��Z��Z�?�x����?7�C!���??!��O��?`��;�?|a���?a���{�?��+Q��?�]�ڕ��?              �?      �?      �?              �?۶m۶m�?I�$I�$�?      �?      �?      �?      �?      �?                      �?      �?                      �?ZZZZZZ�?�������?9��8���?�q�q�?      �?      �?      �?        333333�?�������?              �?      �?              �?                      �?�������?�������?eMYS֔�?MYS֔5�?      �?      �?(������?6��P^C�?      �?      �?              �?�$I�$I�?۶m۶m�?              �?      �?                      �?�������?�������?;�;��?�؉�؉�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?333333�?�������?ffffff�?              �?(�����?�5��P�?�$I�$I�?۶m۶m�?      �?                      �?              �?DDDDDD�?wwwwww�?333333�?�������?              �?      �?        ffffff�?333333�?�$I�$I�?۶m۶m�?      �?        �������?333333�?      �?      �?              �?      �?                      �?      �?        �������?�������?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?4u~�!��?Y1P�M�?      �?        ��+Q��?�]�ڕ��?              �?^Cy�5�?(������?�q�q�?�q�q�?(������?6��P^C�?      �?      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?        AZ��@�?���o)��?:����?���=��?o���o�?�r�!��?�}��?��Gp�?�m۶m��?�$I�$I�?              �?ى�؉��?�؉�؉�?      �?      �?�m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?                      �?      �?        qG�w��?w�qGܱ?�������?�?      �?      �?      �?      �?      �?                      �?      �?              �?        ;�;��?;�;��?      �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        :�h�́�?2~�ԓ�?      �?      �?#�u�)��?v�)�Y7�?UUUUUU�?UUUUUU�?              �?      �?        KKKKKK�?�������?      �?              �?      �?;�;��?ى�؉��?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?n۶m۶�?�$I�$I�?O��N���?;�;��?      �?        ffffff�?�������?��8��8�?�q�q�?n۶m۶�?�$I�$I�?      �?              �?              �?      �?              �?      �?        ��sH�?�琚`��?uo@����?[��5;j�?      �?        w�qG�?qG�wĽ?      �?      �?      �?      �?[k���Z�?�RJ)���?(������?^Cy�5�?      �?              �?      �?              �?      �?        ⎸#��?w�qG��?333333�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?        >����?|���?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?              �?      �?              �?        �����? �����?�������?�?/�袋.�?F]t�E�?      �?        xxxxxx�?�?      �?      �?              �?      �?        ;�;��?;�;��?      �?              �?      �?      �?        |�W|�W�?�A�A�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?�������?333333�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?        Lg1��t�?g1��t�?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?        ��O��O�?l�l��?      �?        >���>�?|���?�������?333333�?�$I�$I�?۶m۶m�?              �?�������?�������?      �?      �?      �?                      �?      �?                      �?ӛ���7�?d!Y�B�?      �?        �������?�������?333333�?�������?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ��sHM�?:�&oe�?              �?���
b�?m�w6�;�?�������?�?�������?�?      �?      �?              �?ى�؉��?�؉�؉�?      �?      �?      �?      �?      �?                      �?      �?        333333�?�������?              �?      �?      �?      �?                      �?�������?333333�?      �?              �?      �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?                      �?      �?        vb'vb'�?;�;��?      �?      �?�������?�������?              �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���bhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       j                    �?v�_���?�           8�@               i                 p�H@�+����?�            �k@              `                 0C�>@����)��?n            �e@                                 �1@�xO��(�?b             c@                                ���,@$�q-�?             :@        ������������������������       �                     &@                                   �?�r����?
             .@              	                     @�C��2(�?             &@        ������������������������       �                     @        
                           �?      �?             @                               `�@1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?               S                 Ь�9@PlX=��?Q            �_@              .                   �;@
j*D>�?B             Z@               '                   �6@b�2�tk�?             B@                                 �2@�G��l��?             5@                                   �?      �?              @                               P��@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                  �3@�	j*D�?	             *@        ������������������������       �                      @                                   �?���|���?             &@        ������������������������       �                      @                                   �4@X�<ݚ�?             "@        ������������������������       �                     �?        !       $                   �5@      �?              @        "       #                 03S$@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        %       &                 �̜!@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        (       )                 ��Y#@z�G�z�?	             .@        ������������������������       �                     @        *       +                 0S�-@      �?              @        ������������������������       �                      @        ,       -                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        /       4                    �?�!���?,             Q@        0       1                 �%@      �?              @        ������������������������       �                     �?        2       3                 �|Y=@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        5       >                     @��0u���?&             N@        6       =                    �?�����?             5@       7       8                    �?�����H�?	             2@        ������������������������       �                      @        9       <                 `f&'@      �?             0@        :       ;                   �J@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        ?       D                    �?�n_Y�K�?            �C@       @       A                 ���@R���Q�?             4@        ������������������������       �                      @        B       C                    �?�X�<ݺ?             2@       ������������������������       �                     1@        ������������������������       �                     �?        E       P                    @@p�ݯ��?             3@       F       G                 �|�<@����X�?	             ,@        ������������������������       �                      @        H       M                 �|Y>@�q�q�?             (@       I       L                 pf�3@      �?              @       J       K                 pf&(@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        N       O                 03C3@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        Q       R                   @B@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        T       [                 ��9;@�㙢�c�?             7@       U       V                   @C@�X�<ݺ?             2@       ������������������������       �                     &@        W       X                     �?؇���X�?             @        ������������������������       �                     @        Y       Z                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        \       _                     @���Q��?             @        ]       ^                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        a       b                     @����X�?             5@        ������������������������       �                     @        c       d                 ��T?@�t����?             1@        ������������������������       �                      @        e       h                    @�<ݚ�?             "@       f       g                 ��p@@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        #             H@        k       �                    �?��]��?6           �~@       l       �                     �?T�6|���?            z@        m       ~                    �?�)
;&��?6             W@        n       }                 p�w@���Q��?             >@       o       |                 @�pX@X�Cc�?             <@       p       {                   @J@�q�q�?             8@       q       z                    C@X�<ݚ�?             2@       r       w                  Y>@և���X�?	             ,@       s       v                 ���<@      �?              @       t       u                 ��";@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        x       y                 @�6M@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @               �                 03�U@�&�5y�?#             O@       �       �                   @L@>���Rp�?              M@       �       �                   �>@�q�q�?             H@        �       �                   �9@
;&����?             7@        ������������������������       �                     @        �       �                   �=@      �?             0@       �       �                 `f�;@�q�q�?             (@       �       �                   @G@z�G�z�?             $@       �       �                 03k:@����X�?             @        ������������������������       �                      @        ������������������������       ����Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @B@HP�s��?             9@       ������������������������       �        	             (@        �       �                   �E@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     $@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���x&�?�            @t@        �       �                 �y�'@4?,R��?.             R@       �       �                 pF�#@r�q��?"             K@       �       �                    �?f1r��g�?!            �J@       �       �                   @@6YE�t�?            �@@       �       �                   �6@��s����?             5@        ������������������������       �                      @        �       �                 ���@�KM�]�?             3@       ������������������������       �                     &@        �       �                 �|=@      �?              @        ������������������������       �                      @        �       �                 �|�=@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        �       �                 �|Y=@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                  ��@R���Q�?             4@        ������������������������       �                     "@        �       �                 �|Y=@���!pc�?	             &@        ������������������������       �                      @        �       �                 X��A@�����H�?             "@       ������������������������       �؇���X�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     @�X�<ݺ?             2@        ������������������������       �                     @        �       �                    �?�8��8��?             (@        ������������������������       �                     @        �       �                   `3@z�G�z�?             @        ������������������������       �                      @        �       �                 03�7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @@@�8��8��?�            �o@       �       �                     @ .2��A�?x            �g@        �       �                 �|Y=@     ��?             @@       ������������������������       �                     2@        �       �                 �|�=@d}h���?             ,@        �       �                    @      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �>@��-�=��?`            �c@       �       �                 �?�@Hm_!'1�?Z            `b@       �       �                 �?$@P�Lt�<�?/             S@        �       �                    7@�7��?            �C@       ������������������������       �                     :@        �       �                 ���@8�Z$���?
             *@        �       �                 �&b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���@ףp=
�?             $@       ������������������������       �                     @        �       �                 �|�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �B@        �       �                 �|Y=@D��\��?+            �Q@       �       �                   �:@��<b���?             G@       �       �                   �3@�?�'�@�?             C@        �       �                 ��Y @�	j*D�?	             *@        �       �                   �2@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                      @        �       �                   �4@`2U0*��?             9@        �       �                 @3�@      �?              @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     1@        �       �                   �;@      �?              @        ������������������������       �                     @        �       �                 �̌!@���Q��?             @        ������������������������       �                      @        �       �                   �<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     9@        �       �                 �!B@X�<ݚ�?             "@       �       �                 �?�@����X�?             @        ������������������������       �                      @        �       �                 pf�'@���Q��?             @       �       �                   �?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                     @      �?)             P@        �       �                    1@ 7���B�?             ;@       �       �                 `f�)@      �?
             0@        ������������������������       �                     @        �       �                   @D@ףp=
�?             $@        ������������������������       �                     @        �       �                   �F@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                 �?�@�?�|�?            �B@       ������������������������       �                     9@        �       �                 @3�@�8��8��?
             (@        ������������������������       �      �?              @        ������������������������       �                     $@        �                       @3�4@z�7�Z�?1            @R@        �       �                     @���!pc�?             6@        ������������������������       �                     @                               H�^ @�q�q�?             2@        ������������������������       �                      @                                 �?      �?             0@        ������������������������       �                      @                                �*@����X�?	             ,@        ������������������������       �                     @                                �1@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        	                         �?��x_F-�?#            �I@        
                         8@�q�q�?	             .@        ������������������������       �                     @                              tՌs@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?                                 �?4?,R��?             B@        ������������������������       �                     @                                 @     ��?             @@                                  @�q�q�?	             (@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     4@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������ *�3�?���M���?�+c���?jNq��?[�~�u��?R�@&��?�?�?��?6��5���?;�;��?�؉�؉�?              �?�?�������?F]t�E�?]t�E�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?        ��`0�?�|>����?;�;��?b'vb'v�?�8��8��?9��8���?��y��y�?1�0��?      �?      �?      �?      �?              �?      �?              �?        ;�;��?vb'vb'�?              �?F]t�E�?]t�E]�?              �?�q�q�?r�q��?      �?              �?      �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?              �?      �?              �?�������?UUUUUU�?              �?      �?        �������?�������?      �?      �?              �?�m۶m��?�$I�$I�?              �?      �?        """"""�?�������?�a�a�?=��<���?�q�q�?�q�q�?              �?      �?      �?�$I�$I�?�m۶m��?              �?      �?                      �?              �?ى�؉��?;�;��?333333�?333333�?      �?        �q�q�?��8��8�?              �?      �?        ^Cy�5�?Cy�5��?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?�������?333333�?      �?                      �?      �?              �?      �?      �?                      �?�������?333333�?              �?      �?        d!Y�B�?�7��Mo�?�q�q�?��8��8�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �m۶m��?�$I�$I�?              �?<<<<<<�?�?      �?        9��8���?�q�q�?�m۶m��?�$I�$I�?              �?      �?              �?                      �?8͸G_�?����?'vb'vb�?b'vb'v�?���7���?C���,�?333333�?�������?%I�$I��?�m۶m��?�������?�������?�q�q�?r�q��?�$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?                      �?�������?UUUUUU�?      �?                      �?              �?      �?              �?                      �?:�s�9�?�1�c��?�i��F�?GX�i���?�������?�������?�Mozӛ�?Y�B��?      �?              �?      �?UUUUUU�?UUUUUU�?�������?�������?�$I�$I�?�m۶m��?              �?�������?333333�?              �?      �?                      �?q=
ףp�?{�G�z�?      �?        ;�;��?;�;��?              �?      �?              �?              �?      �?      �?                      �?��a�2��?�2�tk~�?�8��8��?r�q��?�������?UUUUUU�?�!5�x+�?�x+�R�?'�l��&�?e�M6�d�?z��y���?�a�a�?              �?�k(���?(�����?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        333333�?333333�?      �?        F]t�E�?t�E]t�?              �?�q�q�?�q�q�?۶m۶m�?�$I�$I�?      �?                      �?��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?�+����?g���Q߹?      �?      �?      �?        I�$I�$�?۶m۶m�?      �?      �?      �?                      �?      �?        }˷|˷�?�A�A�?Y�Cc�?9/���?���k(�?(�����?��[��[�?�A�A�?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �o�z2~�?�@�6�?��,d!�?��Moz��?������?y�5���?vb'vb'�?;�;��?�������?�������?              �?UUUUUU�?UUUUUU�?      �?        ���Q��?{�G�z�?      �?      �?      �?      �?      �?              �?              �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        r�q��?�q�q�?�m۶m��?�$I�$I�?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?	�%����?h/�����?      �?      �?      �?        �������?�������?      �?        �������?�������?              �?      �?              �?        *�Y7�"�?к����?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        �I�&M��?�lٲe��?t�E]t�?F]t�E�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?�$I�$I�?�m۶m��?              �?F]t�E�?]t�E]�?              �?      �?        �������?�?UUUUUU�?UUUUUU�?              �?]t�E�?F]t�E�?      �?                      �?�8��8��?r�q��?      �?              �?      �?�������?�������?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ+�MhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0Kh2h3h4hph<�h=Kub��������       T                    �?�s�ˈ.�?�           8�@                                    @衶� �?�            @o@              
                     �?���?Z            �`@                                  "@P�Lt�<�?/             S@        ������������������������       �                     �?               	                 �DD@�}��L�?.            �R@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        )            �P@                                  �*@�j��b�?+            �M@                                  �J@��s����?             5@                               ��Y)@�KM�]�?             3@        ������������������������       �                     $@                                   5@�<ݚ�?             "@        ������������������������       �                      @                                   :@����X�?             @        ������������������������       �                     �?                                   B@r�q��?             @       ������������������������       �                     @                                   D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                  �E@�}�+r��?             C@       ������������������������       �                     >@                                  �8@      �?              @        ������������������������       �                     @                                  @F@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                '                    �?
;&����?E            �\@        !       &                 X�,A@4?,R��?             B@       "       #                    �?l��\��?             A@       ������������������������       �                     =@        $       %                 �|Y=@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        (       G                 ���1@t�C�#��?.            �S@       )       B                 ��Y.@Tt�ó��?            �H@       *       ?                    �?�s��:��?             C@       +       .                 pf�@և���X�?             <@        ,       -                 �|Y:@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        /       8                   �9@      �?             6@       0       3                   �3@�q�q�?	             (@        1       2                 �&B@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        4       5                   �5@      �?              @        ������������������������       �                     @        6       7                   �6@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        9       >                   �C@�z�G��?             $@       :       ;                 @3�@      �?              @        ������������������������       �                     @        <       =                 �|�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        @       A                    7@      �?             $@       ������������������������       �                     @        ������������������������       �                     @        C       F                 �|�;@�C��2(�?             &@        D       E                 pff0@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        H       M                    �?��S�ۿ?             >@        I       J                    �?      �?              @        ������������������������       �                     @        K       L                 ���4@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        N       S                 ��p@@���7�?             6@       O       P                   �8@�����H�?             "@       ������������������������       �                     @        Q       R                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        U       �                     �?O��,4�?'           �|@        V       m                  �>@�I� �?:             W@        W       ^                    �?|��?���?             ;@        X       Y                 �|�=@      �?             @        ������������������������       �                     �?        Z       [                   @@@�q�q�?             @        ������������������������       �                     �?        \       ]                    <@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        _       f                   �@@
;&����?             7@        `       a                   �<@z�G�z�?             $@        ������������������������       �                     �?        b       c                 `fF<@�����H�?             "@       ������������������������       �                     @        d       e                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        g       l                   �H@�θ�?	             *@       h       i                   �9@      �?              @        ������������������������       �                      @        j       k                    D@r�q��?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     @        n       �                 �̾w@؇>���?&            @P@       o       v                    �?     ��?%             P@        p       s                  �}S@      �?             @@        q       r                   @J@      �?             $@       ������������������������       �                     @        ������������������������       �                     @        t       u                   �1@��2(&�?	             6@        ������������������������       �                     @        ������������������������       �                     3@        w       x                    �?     ��?             @@        ������������������������       �                     �?        y       �                 03�T@��a�n`�?             ?@       z       �                    F@8�Z$���?             :@       {       �                  x#J@      �?
             0@       |                        ��yC@ףp=
�?             $@        }       ~                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �C@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                 ~�.@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                 �w|c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @4Qi0���?�            w@        �       �                    "@`-�I�w�?1             S@        ������������������������       �                     �?        �       �                 �|Y=@Х-��ٹ?0            �R@        ������������������������       �                     7@        �       �                    �?$�q-�?!             J@       �       �                 �|�=@HP�s��?             I@        �       �                    @�<ݚ�?             "@       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @D@������?            �D@        ������������������������       �                     5@        �       �                   �*@ףp=
�?             4@        �       �                 `f�)@"pc�
�?             &@        ������������������������       �                     @        �       �                   �F@�q�q�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        �       �                 ��) @��T �?�            Pr@       �       �                    �?8��$��?w            �g@        �       �                    �?���5��?#            �L@       �       �                 �|Y=@$G$n��?            �B@        �       �                   @@�q�q�?             .@       �       �                    �?�θ�?             *@       �       �                 ��y@      �?             (@        ������������������������       �                     @        �       �                   �6@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        �       �                 X��A@ףp=
�?             4@       �       �                 ���@�t����?             1@        ������������������������       �                     @        �       �                 ��(@8�Z$���?
             *@       ������������������������       �r�q��?	             (@        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@�\=lf�?T            �`@       �       �                    �?�ջ����?@             Z@       �       �                 ���@@�n���??            �Y@        �       �                   �8@Pa�	�?            �@@        �       �                 ���@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �        .            �Q@        ������������������������       �                     �?        �       �                 @3�@(;L]n�?             >@        �       �                   �4@�C��2(�?             &@        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     3@        �       �                    �?�4�M�f�?E            �Y@       �       �                    �?��!���??            @W@       �       �                    �?@�0�!��?-             Q@        �       �                   �:@�q�q�?             (@        �       �                    '@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 0SE @؇���X�?&             L@        ������������������������       �                     �?        �       �                   �9@X�;�^o�?%            �K@        ������������������������       �                     4@        �       �                   �;@z�G�z�?            �A@        ������������������������       �                     @        �       �                 �|�=@��a�n`�?             ?@       �       �                    (@���N8�?             5@        �       �                   �<@z�G�z�?             @        ������������������������       �                     �?        �       �                 �|Y=@      �?             @       �       �                 ���"@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             0@        �       �                 �T)D@z�G�z�?             $@       �       �                 ��)"@�����H�?             "@        ������������������������       �                     @        �       �                 ���'@z�G�z�?             @        �       �                   �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    0@ �o_��?             9@        �       �                 `ff/@�<ݚ�?             "@       �       �                 �|�?@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     0@        ������������������������       �                     "@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub���������������0Ȍ��?��o��?T㥛� �?V-����?t��:W�?��oS��?(�����?���k(�?      �?        O贁N�?�_,�Œ�?      �?      �?      �?                      �?              �?��/���?�N��?�a�a�?z��y���?(�����?�k(���?              �?�q�q�?9��8���?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        (�����?�5��P�?              �?      �?      �?              �?�������?333333�?      �?                      �?�Mozӛ�?Y�B��?r�q��?�8��8��?�������?------�?              �?333333�?�������?              �?      �?              �?        ��td�@�?��7a~�?/�����?h�����?��k(��?�k(���?�$I�$I�?۶m۶m�?�������?UUUUUU�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?        333333�?ffffff�?      �?      �?              �?      �?      �?      �?                      �?      �?              �?      �?              �?      �?        F]t�E�?]t�E�?      �?      �?      �?                      �?              �?�������?�?      �?      �?      �?              �?      �?              �?      �?        �.�袋�?F]t�E�?�q�q�?�q�q�?      �?              �?      �?      �?                      �?      �?        ���c|��?�l,p~�?Y�B���?Nozӛ��?	�%����?{	�%���?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �Mozӛ�?Y�B��?�������?�������?              �?�q�q�?�q�q�?      �?              �?      �?      �?                      �?�؉�؉�?ى�؉��?      �?      �?      �?        UUUUUU�?�������?              �?      �?      �?              �?�����? �����?     ��?      �?      �?      �?      �?      �?              �?      �?        ��.���?t�E]t�?              �?      �?              �?      �?      �?        �c�1��?�s�9��?;�;��?;�;��?      �?      �?�������?�������?      �?      �?      �?                      �?      �?              �?      �?      �?                      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?#6�a#�?�On��?Q^Cy��?y�5�װ?              �?K~��K�?O贁N�?      �?        �؉�؉�?;�;��?q=
ףp�?{�G�z�?9��8���?�q�q�?      �?              �?      �?      �?                      �?p>�cp�?������?      �?        �������?�������?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?              �?        �H�%��?ڻ�p�v�?vX�Q�}�?�x��* �?�}��?��Gp�?к����?���L�?UUUUUU�?UUUUUU�?ى�؉��?�؉�؉�?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?                      �?      �?        �������?�������?<<<<<<�?�?      �?        ;�;��?;�;��?�������?UUUUUU�?      �?              �?        "=P9���?g��1��?;�;��?;�;��?\mMw��?��,�?|���?|���?�؉�؉�?;�;��?      �?                      �?      �?              �?              �?        �������?�?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?              �?        





�?�������?v�e�]v�?'�h��&�?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?      �?        ۶m۶m�?�$I�$I�?              �?�־a��?J��yJ�?      �?        �������?�������?              �?�s�9��?�c�1Ƹ?��y��y�?�a�a�?�������?�������?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?�q�q�?�q�q�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?
ףp=
�?�Q����?�q�q�?9��8���?�������?333333�?              �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJY]hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       4                     �?�����?�           8�@                                   �?���}��?b             c@        ������������������������       �        +            @Q@               1                    �?��q7L��?7            �T@              ,                    K@ꮃG��?.            @Q@                                 �9@�p����?)            �N@        ������������������������       �                     @                                 �>@��>4և�?%             L@        	                        ���<@؇���X�?             5@       
                           �?�z�G��?             $@        ������������������������       �                     �?                                03k:@�<ݚ�?             "@        ������������������������       �                      @                                �|�?@����X�?             @                                �|�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �C@z�G�z�?             @        ������������������������       �                      @                                  @G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     &@               '                    H@�xGZ���?            �A@                                 �;@�q�q�?             ;@                                   6@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                                  @K@      �?             4@       ������������������������       �        	             &@               "                    �?X�<ݚ�?             "@                !                 p�w@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        #       $                 03�M@�q�q�?             @        ������������������������       �                      @        %       &                 03�U@      �?             @       ������������������������       �                      @        ������������������������       �                      @        (       )                   �H@      �?              @        ������������������������       �                     @        *       +                 ���W@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        -       .                 ���=@      �?              @        ������������������������       �                     @        /       0                   �R@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        2       3                   @B@X�Cc�?	             ,@        ������������������������       �                     @        ������������������������       �                     "@        5       r                    �?�9����?j           x�@        6       C                   �6@��+��?Y            �b@        7       @                  18@���B���?             :@       8       9                 P��+@�}�+r��?             3@       ������������������������       �                     *@        :       ?                    �?r�q��?             @       ;       <                   �@z�G�z�?             @        ������������������������       �                      @        =       >                   �-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        A       B                     @և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        D       M                 ���@6}��#�?H            �^@        E       F                 ���@XB���?             =@       ������������������������       �        
             ,@        G       H                 �|=@��S�ۿ?	             .@        ������������������������       �                     @        I       L                 ���@ףp=
�?             $@       J       K                 �|�=@؇���X�?             @       ������������������������       �r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        N       q                 `v�9@��MΖ��?5            @W@       O       p                    �?��9܂�?1            @V@       P       m                    �?�)��V��?/            �T@       Q       V                    �?D�n�3�?+             S@        R       S                   @,@Pa�	�?            �@@       ������������������������       �                     5@        T       U                  S�-@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        W       b                 �|Y=@^����?            �E@        X       _                    �?      �?             (@       Y       Z                     @      �?             $@        ������������������������       �                     @        [       ^                    <@����X�?             @       \       ]                 �0@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        `       a                  ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        c       l                 �|�=@�n`���?             ?@       d       e                    �?      �?             8@        ������������������������       �                      @        f       k                   `3@���!pc�?             6@       g       j                   @'@z�G�z�?
             4@       h       i                 ���@      �?             0@        ������������������������       �                     �?        ������������������������       �������?             .@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        n       o                 03�-@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        s       �                    �?�����?           �y@        t       �                 ���P@8��~P�?P            �^@       u       z                    !@�m���?N            �]@        v       w                 03�<@�}�+r��?             3@       ������������������������       �                     &@        x       y                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        {       �                 03�;@4���C�?B            �X@       |       �                    :@Pi�����?9            �T@       }       �                   �>@���L��?5            �S@       ~                          �1@~|z����?"            �J@        ������������������������       �                     @        �       �                     @�`���?             �H@        �       �                    �?�<ݚ�?             "@       �       �                   �;@���Q��?             @       �       �                   �6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?H�z�G�?             D@       �       �                   �@l��[B��?             =@        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 Ь�#@�q�q�?             5@        ������������������������       �                      @        �       �                 03�0@��
ц��?             *@       �       �                 �|�9@      �?              @        �       �                 �[$@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �;@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        �       �                     @�+e�X�?             9@       �       �                    L@�<ݚ�?             2@       �       �                   �B@      �?             0@       ������������������������       �                     $@        �       �                    D@�q�q�?             @        ������������������������       �                     �?        �       �                    5@z�G�z�?             @       ������������������������       �                     @        �       �                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ��Y.@����X�?             @       �       �                  SE"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                     @     ��?	             0@        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        �       �                    @�%��5�?�            r@        �       �                   �C@      �?             0@       �       �                    �?؇���X�?	             ,@       �       �                    @�C��2(�?             &@       �       �                 ���7@r�q��?             @        �       �                 �(\�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �T�I@($�pa�?�            q@       �       �                 P�N@X�l�ؾ?�            �p@        ������������������������       �        *             L@        �       �                     @,�T�6�?�             j@        �       �                    @@��GEI_�?&            �N@        ������������������������       �                     6@        �       �                    �?��-�=��?            �C@       �       �                    F@      �?             @@        �       �                   �3@����X�?	             ,@       �       �                   �'@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   @D@      �?              @       �       �                   @B@z�G�z�?             @       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                     @        �       �                    �?�1h�'��?_            `b@       �       �                 �Yu@��ׄ��?Z            `a@        �       �                    �?�q�q�?             @       �       �                    =@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    '@���D�k�?W            �`@        �       �                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?0�v���?U            ``@       �       �                   �0@6uH���?O             _@        �       �                 �̌!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �:@\����?L            @^@        ������������������������       �                     @@        �       �                   �;@ą%�E�?5            @V@        ������������������������       �                      @        �       �                 �|�=@����?4            �U@       �       �                   �<@0G���ջ?             J@        ������������������������       �                     @        �       �                 �|Y=@��S�ۿ?            �F@        �       �                 ���"@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��) @@-�_ .�?            �B@       ������������������������       �                     8@        �       �                 pf� @8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        �       �                 @3�@(N:!���?            �A@        �       �                 �?�@z�G�z�?
             .@        ������������������������       �                     "@        �       �                   �?@      �?             @        ������������������������       �                     �?        �       �                   �A@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �      �?              @        �       �                   �"@P���Q�?             4@       ������������������������       �        	             ,@        �       �                    ?@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �                            @�q�q�?             "@        ������������������������       �                     �?                                 ;@      �?              @        ������������������������       �                      @                              p�O@r�q��?             @                             �|�>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������w��	�?�3����?������?(������?              �?��\V��?��FS���?�%~F��?s��\;�?C��6�S�?ާ�d��?      �?        I�$I�$�?۶m۶m�?�$I�$I�?۶m۶m�?333333�?ffffff�?      �?        �q�q�?9��8���?              �?�$I�$I�?�m۶m��?      �?      �?              �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?              �?              �?�_�_�?�A�A�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?      �?      �?      �?        �q�q�?r�q��?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?%I�$I��?�m۶m��?              �?      �?        � �*���?��Ѫe~�?�S�n�?*�Y7�"�?ى�؉��?��؉���?(�����?�5��P�?              �?UUUUUU�?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?۶m۶m�?              �?      �?        �u�y��?�����?GX�i���?�{a���?      �?        �������?�?      �?        �������?�������?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?              �?        �]v�e��?4�DM4�?�.p��? ��G?��?GS��r�?]V��F�?(������?l(�����?|���?|���?              �?UUUUUU�?UUUUUU�?      �?                      �?�qG��?w�qG��?      �?      �?      �?      �?      �?        �$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?�9�s��?�c�1��?      �?      �?      �?        F]t�E�?t�E]t�?�������?�������?      �?      �?      �?        wwwwww�?�?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?              �?        ؿ$J��?P���k��?�`mާ�?�Oq���?ylE�pR�?�Iݗ�V�?(�����?�5��P�?              �?      �?      �?      �?                      �?'�l��&�?m��&�l�?��FS��?���\V�?��o��o�?�4H�4H�?��sHM0�?�	�[���?              �?����S�?և���X�?�q�q�?9��8���?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?ffffff�?333333�?���=��?GX�i���?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?        �؉�؉�?�;�;�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        F]t�E�?t�E]t�?              �?      �?        ���Q��?R���Q�?�q�q�?9��8���?      �?      �?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?              �?      �?              �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?              �?      �?              �?        �V�e�t�?�IєX�?      �?      �?�$I�$I�?۶m۶m�?F]t�E�?]t�E�?UUUUUU�?�������?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        ~ڧ}ڧ�?,�,��?��|��?|��|�?      �?        'vb'vb�?�N��N�?�d����?;ڼOqɰ?      �?        }˷|˷�?�A�A�?      �?      �?�m۶m��?�$I�$I�?r�q��?�q�q�?      �?              �?      �?�������?�������?      �?      �?      �?                      �?      �?              �?              �?        K���+�?�E�_���?�Ke{��?��$D�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �՝VwZ�?�RKE,�?      �?      �?      �?                      �?�2����?�i��?k���Zk�?��RJ)��?UUUUUU�?UUUUUU�?              �?      �?        ���|���?"pc�
�?      �?        �as���?��g<�?              �?��֡�l�?/�I���?vb'vb'�?�؉�؉�?      �?        �������?�?      �?      �?      �?                      �?S�n0E�?к����?      �?        ;�;��?;�;��?              �?      �?        |�W|�W�?�A�A�?�������?�������?      �?              �?      �?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?ffffff�?�������?      �?        �������?UUUUUU�?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ4
hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������                           @��eC~�?�           8�@                                   �?���!pc�?            �@@        ������������������������       �                     @                                   �?8^s]e�?             =@                                  �?z�G�z�?             4@                                   @ףp=
�?             $@        ������������������������       �                     @               	                     @z�G�z�?             @        ������������������������       �                      @        
                           �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                    @�z�G��?             $@        ������������������������       �                     @                                ��|2@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                   �?X�<ݚ�?             "@                                   @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                �Q��?�q�q�?             @        ������������������������       �                     �?                                pf�C@z�G�z�?             @                                  @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               �                     @���P���?�           0�@               e                 ���=@\������?�             t@              >                    �?�&!��?l            �e@                #                     �?6YE�t�?'            �P@        !       "                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        $       1                   �*@     ��?%             P@        %       (                 ��Y)@     ��?             @@       &       '                   �J@�KM�]�?	             3@       ������������������������       �                     1@        ������������������������       �                      @        )       ,                    <@�	j*D�?             *@        *       +                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        -       .                   �B@�����H�?             "@       ������������������������       �                     @        /       0                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        2       =                    �?     ��?             @@       3       4                   �2@      �?             8@        ������������������������       �                     @        5       8                   �6@@�0�!��?             1@        6       7                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        9       :                    9@؇���X�?	             ,@        ������������������������       �                     �?        ;       <                   �E@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                      @        ?       d                    �?���C��?E            �Z@       @       W                 ��$:@      �??             X@       A       B                     �?`2U0*��?3            �R@        ������������������������       �                     @        C       D                    �?hA� �?/            �Q@        ������������������������       �                     @        E       J                    5@     �?+             P@        F       G                   �2@r�q��?             @        ������������������������       �                      @        H       I                   �'@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        K       V                   �E@XB���?&             M@       L       M                   �'@���N8�?             E@        ������������������������       �                     0@        N       U                   @D@$�q-�?             :@       O       T                 �|�=@ �q�q�?             8@        P       S                    1@�����H�?             "@       Q       R                 �|�<@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             .@        ������������������������       �      �?              @        ������������������������       �                     0@        X       c                 `f�:@և���X�?             5@       Y       Z                    �?�	j*D�?             *@        ������������������������       �                     �?        [       \                 03k:@�q�q�?             (@        ������������������������       �                     @        ]       ^                   �C@X�<ݚ�?             "@        ������������������������       �                     @        _       `                   @G@�q�q�?             @        ������������������������       �                      @        a       b                    K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        f       �                    @�y��?�?[            �b@       g       h                  �>@���X��?Z            �b@        ������������������������       �                     ,@        i       j                    �?R��	P�?T            �`@        ������������������������       �        *            �O@        k       �                     �?�E��ӭ�?*             R@       l       s                  x#J@:ɨ��?&            �P@        m       n                    �?�LQ�1	�?             7@        ������������������������       �                     @        o       r                 ��yC@@�0�!��?	             1@        p       q                   @A@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        t       �                 Ј@S@�&!��?            �E@        u       ~                    F@�û��|�?             7@       v       w                    5@؇���X�?             ,@        ������������������������       �                     �?        x       }                 `f�K@$�q-�?             *@        y       z                 `�iJ@r�q��?             @        ������������������������       �                     @        {       |                    @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               �                   �H@�<ݚ�?             "@        �       �                   �G@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?R���Q�?             4@       �       �                 �̾w@�����H�?
             2@       �       �                 ���X@�IєX�?	             1@        �       �                    ?@z�G�z�?             @        ������������������������       �                      @        �       �                    G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     �?        �       �                    6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��0�]��?�            @v@        �       �                   �-@�����?A            �Z@        ������������������������       �                     *@        �       �                    �?      �?:            �W@       �       �                    �?h+�v:�?)             Q@        �       �                    �?6YE�t�?            �@@        �       �                 �|Y6@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���@ �Cc}�?             <@        ������������������������       �                     @        ������������������������       �                     9@        �       �                   �@���Q��?            �A@        �       �                    8@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                  �#@l��
I��?             ;@        �       �                   �9@@4և���?             ,@       ������������������������       �                     $@        �       �                    ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�;@��
ц��?	             *@       �       �                 �[$@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��1@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @C@���B���?             :@       �       �                 ���5@�t����?             1@        �       �                   �/@���Q��?             @       �       �                    �?�q�q�?             @       �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 pVm<@r�q��?             (@        ������������������������       �                     @        �       �                 X��@@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        �       �                   @@@�cX1!��?�             o@       �       �                   �?@ i���t�?�            �h@       �       �                    �?�! �	��?�            �g@        �       �                    �?p�ݯ��?             3@       �       �                   �5@؇���X�?             ,@        ������������������������       �                      @        ������������������������       �        
             (@        ������������������������       �                     @        �       �                 �|�=@���@�c�?r            �e@       �       �                   �:@�ۊ�̴?o            �d@       �       �                   @4@�|���?<             V@        �       �                    �?@��8��?             H@       �       �                   �3@(;L]n�?             >@       ������������������������       �                     2@        �       �                 @3�@�8��8��?	             (@       �       �                 P�@z�G�z�?             @       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        	             2@        ������������������������       �                     D@        �       �                 �?$@�S(��d�?3            @S@        �       �                    �?�㙢�c�?             7@       �       �                  s�@     ��?
             0@        ������������������������       �                     @        �       �                 �|Y=@���!pc�?             &@        ������������������������       �                     �?        ������������������������       �z�G�z�?             $@        �       �                 ��@؇���X�?             @       ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                   �;@ 7���B�?$             K@        �       �                 �� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �? pƵHP�?"             J@       �       �                 ���"@p���?              I@       ������������������������       �                     C@        �       �                 �|Y=@�8��8��?
             (@        �       �                   �<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        �       �                 �̌!@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 P�@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                    �J@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub����������������Kkz�?�fh)�?t�E]t�?F]t�E�?              �?	�=����?|a���?�������?�������?�������?�������?              �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        333333�?ffffff�?              �?333333�?�������?              �?      �?        r�q��?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?              �?      �?              �?        g�Pw��?1e^S��?<�?�x4�?�2���e�?֔5eMY�?S֔5eM�?e�M6�d�?'�l��&�?      �?      �?      �?                      �?      �?     ��?      �?      �?(�����?�k(���?              �?      �?        ;�;��?vb'vb'�?      �?      �?      �?                      �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?              �?�������?ZZZZZZ�?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?;�;��?;�;��?              �?      �?                      �?\�琚`�?"5�x+��?      �?      �?���Q��?{�G�z�?      �?        ���?_�_�?      �?             ��?      �?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?        GX�i���?�{a���?��y��y�?�a�a�?      �?        �؉�؉�?;�;��?�������?UUUUUU�?�q�q�?�q�q�?�������?�������?      �?                      �?      �?              �?              �?      �?      �?        �$I�$I�?۶m۶m�?;�;��?vb'vb'�?              �?UUUUUU�?UUUUUU�?              �?�q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?        �6�i��?��K~��?�IA��U�?[���?              �?n�Q�ߦ�?�:W���?              �?�q�q�?r�q��?N6�d�M�?e�M6�d�?��Moz��?Y�B��?      �?        ZZZZZZ�?�������?      �?      �?      �?                      �?      �?        ֔5eMY�?S֔5eM�?��,d!�?8��Moz�?�$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?9��8���?�q�q�?333333�?�������?      �?                      �?      �?        333333�?333333�?�q�q�?�q�q�?�?�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?              �?      �?              �?              �?         ��G?��?�\��?�_����?�@�Ե�?      �?              �?      �?xxxxxx�?�������?e�M6�d�?'�l��&�?�������?333333�?              �?      �?        ۶m۶m�?%I�$I��?      �?                      �?333333�?�������?      �?      �?              �?      �?        Lh/����?h/�����?n۶m۶�?�$I�$I�?      �?              �?      �?              �?      �?        �؉�؉�?�;�;�?�������?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?        ��؉���?ى�؉��?�������?�������?�������?333333�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        I�dn�?��ٌ?/�����?����X�?��uX�Q�?:kP<�q�?^Cy�5�?Cy�5��?۶m۶m�?�$I�$I�?              �?      �?                      �?�5eMYS�?���)kʪ?�^G�u��?��[���?��.���?F]t�E�?UUUUUU�?UUUUUU�?�������?�?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?      �?              �?              �?        ������?��O���?�7��Mo�?d!Y�B�?      �?      �?      �?        F]t�E�?t�E]t�?              �?�������?�������?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?	�%����?h/�����?      �?      �?      �?                      �?'vb'vb�?;�;��?\���(\�?{�G�z�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �m۶m��?�$I�$I�?      �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��;hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K�h2h3h4hph<�h=Kub��������       T                    �?���%&�?�           8�@               G                 �|�=@<��u�?�            �l@                               ��@�q�q�?`             b@                                   �?ףp=
�?             4@              
                 ���@�IєX�?
             1@                                �|Y5@      �?             @        ������������������������       �                      @               	                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@                                �|Y:@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?               <                    �?�4�����?S             _@                                   @\��<�|�?@            �W@                                  6@�&=�w��?!            �J@                                   9@؇���X�?	             ,@        ������������������������       �                      @                                ��m1@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �C@               #                    �?      �?             E@                                   @�θ�?             *@        ������������������������       �                     @                                �&�)@�q�q�?	             "@        ������������������������       �                     @                                  �-@���Q��?             @        ������������������������       �                      @                                 �|Y6@�q�q�?             @        ������������������������       �                     �?        !       "                  S�-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        $       1                   �3@����"�?             =@        %       ,                    �?X�Cc�?
             ,@        &       +                 ��y.@և���X�?             @       '       *                   �2@z�G�z�?             @       (       )                 ��!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        -       .                    @����X�?             @        ������������������������       �                     @        /       0                 @3�2@      �?             @        ������������������������       �                      @        ������������������������       �                      @        2       5                 pff@�r����?
             .@        3       4                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        6       7                    :@$�q-�?             *@        ������������������������       �                     @        8       9                   �&@؇���X�?             @        ������������������������       �                     @        :       ;                 �|Y<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        =       @                     @�f7�z�?             =@        >       ?                    @�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        A       B                 ��Z5@      �?             4@        ������������������������       �                     @        C       D                 ��T?@�t����?
             1@       ������������������������       �                     "@        E       F                 pf�C@      �?              @        ������������������������       �                      @        ������������������������       �                     @        H       I                     @����"$�?7            �U@       ������������������������       �        .            �Q@        J       S                 `f68@��S���?	             .@       K       R                    �?���!pc�?             &@       L       Q                 ���*@      �?              @       M       P                   &@r�q��?             @       N       O                    A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        U       �                     �?\5�+=M�?           ~@        V       �                    �?m#9���?A            @\@       W       �                   @J@      �?;             Z@       X       �                   �G@X�<ݚ�?/            @T@       Y       j                    �?���Q��?*            �Q@        Z       ]                   �8@�+e�X�?             9@        [       \                 ���Q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       i                  �>@؇���X�?             5@        _       h                  Y>@      �?             (@       `       g                    B@"pc�
�?             &@       a       b                 �|�;@ףp=
�?             $@        ������������������������       �                      @        c       f                 �ܵ<@      �?              @       d       e                 X�,@@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        k       �                    �?z�G�z�?            �F@       l       m                 03:@�������?             F@        ������������������������       �                     (@        n       y                   �>@     ��?             @@        o       x                    D@      �?              @       p       w                   @>@����X�?             @       q       v                 `fF<@���Q��?             @       r       s                 03k:@      �?             @        ������������������������       �                     �?        t       u                 �|�<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        z       �                 `f�K@r�q��?             8@       {       |                   �A@�����H�?             2@        ������������������������       �                     @        }       ~                   �B@8�Z$���?	             *@        ������������������������       �                     �?               �                   �;@�8��8��?             (@        �       �                    7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                 03�M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���!pc�?             &@       �       �                 @�pX@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�LQ�1	�?             7@       �       �                   �R@@�0�!��?	             1@       ������������������������       �                     ,@        ������������������������       �                     @        ������������������������       �                     @        �       �                    @�q�q�?             "@       �       �                    6@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @�A����?�             w@        �       �                 �D,C@���Q��?
             .@       �       �                 ���7@"pc�
�?             &@        �       �                 @3�4@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?<{����?�            v@        �       �                 ��� @R���Q�?             D@       �       �                 �|Y=@z�G�z�?             9@        �       �                 ��y@X�<ݚ�?             "@        ������������������������       �                     @        �       �                   @@�q�q�?             @       �       �                 ���@      �?             @        ������������������������       �                     �?        �       �                   �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 ���@      �?
             0@       ������������������������       �                     "@        �       �                   @@؇���X�?             @       �       �                 �|�=@r�q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��S�ۿ?
             .@       ������������������������       �                     (@        �       �                   �6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���q��?�            �s@       �       �                     @�Rl}��?�            Pr@        �       �                 ��Y)@�.ߴ#�?'            �N@        ������������������������       �                     5@        �       �                   �*@��(\���?             D@       �       �                 �|�=@�����H�?             ;@        �       �                 �|Y<@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �        	             *@        �       �                 ���@��Õty�?�             m@        ������������������������       �                     D@        �       �                 0�gE@��8����?q             h@       �       �                    )@�n�Ƌ��?n            `g@        �       �                    �?���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�Ra����?i             f@        �       �                   `3@r�q��?             8@       �       �                   @'@�LQ�1	�?             7@       �       �                 �|Y=@@�0�!��?             1@        ������������������������       �                     @        ������������������������       �        
             ,@        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�KM�]�?[             c@       �       �                   @@@$V�Ap�?V            �a@       �       �                    ?@@1�`�?G            @^@       �       �                 @3�@�S#א��?D            @]@        �       �                 �?$@`Ӹ����?            �F@        �       �                 �|�;@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �C@        �       �                 `�X#@r�q��?*             R@       �       �                 ���"@d}h���?!             L@       �       �                 @3"@Jm_!'1�?            �H@       �       �                 ��) @��k=.��?            �G@       �       �                   �3@     ��?             @@        ������������������������       �                     @        ������������������������       �                     ;@        �       �                   �:@������?             .@       ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                      @        �       �                   �<@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             0@        �       �                 P�@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �                     "@        �       �                 �|�>@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             4@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������g *��?�0���M�?���9E�?�ʇq�.�?�������?�������?�������?�������?�?�?      �?      �?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ��RJ)��?���Zk��?��%N��?��v�@�?�x+�R�?tHM0���?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?�؉�؉�?ى�؉��?              �?UUUUUU�?UUUUUU�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?	�=����?�i��F�?�m۶m��?%I�$I��?۶m۶m�?�$I�$I�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �$I�$I�?�m۶m��?              �?      �?      �?              �?      �?        �������?�?      �?      �?              �?      �?        �؉�؉�?;�;��?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        O#,�4��?a���{�?�q�q�?9��8���?      �?                      �?      �?      �?              �?<<<<<<�?�?      �?              �?      �?              �?      �?        6eMYSִ?YS֔5e�?              �?�������?�?t�E]t�?F]t�E�?      �?      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?        D��z9�?�z9��?04��A�?�ɗ�|�?      �?      �?r�q��?�q�q�?333333�?�������?���Q��?R���Q�?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?F]t�E�?/�袋.�?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?                      �?�������?�������?t�E]t�?/�袋.�?      �?              �?      �?      �?      �?�$I�$I�?�m۶m��?�������?333333�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �������?UUUUUU�?�q�q�?�q�q�?      �?        ;�;��?;�;��?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        t�E]t�?F]t�E�?      �?      �?              �?      �?                      �?��Moz��?Y�B��?ZZZZZZ�?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        C���,�?�Mozӛ�?�������?333333�?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        3����?j.�W�a�?333333�?333333�?�������?�������?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        �������?�?      �?        UUUUUU�?UUUUUU�?              �?      �?        «�.��?�
���?���0��?F�)�V�?�K�`m�?XG��).�?      �?        �������?333333�?�q�q�?�q�q�?      �?      �?      �?                      �?      �?              �?        �FX�i�?��=���?      �?        �������?UUUUUU�?��X͞��?n�ʄm�?]t�E]�?F]t�E�?      �?                      �?]t�E]�?]t�E�?�������?UUUUUU�?��Moz��?Y�B��?ZZZZZZ�?�������?              �?      �?              �?                      �?�k(���?(�����?�#T�ik�?��^���?�X����?���k���?��+��+�?�꡾??�>��?l�l��?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?UUUUUU�?I�$I�$�?۶m۶m�?����X�?������?g���Q��?br1���?      �?      �?              �?      �?        wwwwww�?�?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?              �?      �?              �?      �?              �?              �?        333333�?�������?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJS�)/hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       `                    �?�Wa�O�?�           8�@               !                     @`מ���?�             o@                                 �&@p���?_            �b@                                  �J@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @                                 "�b@hA� �?Y            �a@                                 �B@`J����?L            �^@       	                          �;@�L��ȕ?7            @W@       
                          �:@��<b�ƥ?             G@       ������������������������       �                     F@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �G@                                  @C@ףp=
�?             >@        ������������������������       �                     �?                                �QD@ 	��p�?             =@                                ���;@"pc�
�?	             &@                                ��9@ףp=
�?             $@        ������������������������       �                     @                                   �?r�q��?             @                                 �I@      �?             @                                 �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     2@                                    !@�t����?             1@        ������������������������       �                      @        ������������������������       �                     .@        "       S                 `f:@4��@���?C             Y@       #       0                 �̌@��=A��?4             S@        $       /                    �?�J�4�?             9@       %       .                 X��B@      �?             8@       &       '                    8@���}<S�?             7@        ������������������������       �                     $@        (       )                   �9@8�Z$���?	             *@        ������������������������       �                     �?        *       +                    �?�8��8��?             (@        ������������������������       �                     �?        ,       -                 ���@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        1       <                 `f�%@��.k���?!            �I@        2       9                    �?�����H�?
             2@       3       8                 pf� @$�q-�?             *@        4       5                 �?�@      �?             @        ������������������������       �                     �?        6       7                   �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        :       ;                   �#@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        =       >                   �#@�q�q�?            �@@        ������������������������       �                     "@        ?       J                 �|�;@r�q��?             8@        @       G                 pff0@�<ݚ�?             "@       A       F                    �?؇���X�?             @       B       E                    �?z�G�z�?             @       C       D                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        H       I                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        K       R                    �?������?             .@       L       M                   �>@d}h���?
             ,@       ������������������������       �                     $@        N       Q                    �?      �?             @       O       P                 ���0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        T       W                    @�8��8��?             8@        U       V                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        X       Y                    �?���7�?             6@        ������������������������       �                     �?        Z       [                    @���N8�?             5@       ������������������������       �        	             1@        \       _                 ���A@      �?             @       ]       ^                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        a       �                   �/@J�W�%�?&           �|@       b       c                     @��|C_�?�            �q@        ������������������������       �        %             O@        d       e                 ���@�ͳ ���?�            �k@        ������������������������       �                     8@        f       �                    �?Lvkef�?�            �h@       g       h                 ��@�����H�?}            �g@        ������������������������       �                     @        i       t                 �Y�@��a�n`�?|            @g@        j       m                 ���@������?             1@        k       l                   �7@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        n       o                   �5@����X�?             @        ������������������������       �                     �?        p       q                 �|=@r�q��?             @        ������������������������       �                      @        r       s                 �|�=@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        u       �                 0SE @0u��Fs�?q             e@       v                          �<@8��d�?R             _@        w       ~                   �4@`Ӹ����?!            �F@        x       {                   �3@�<ݚ�?	             "@       y       z                 �?�@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        |       }                 P�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     B@        �       �                    �?p#�����?1            �S@        �       �                 �|Y=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�r����?.            �R@        �       �                 �|Y=@؇���X�?	             ,@        ������������������������       �                      @        ������������������������       �                     (@        �       �                   �D@(��+�?%            �N@       �       �                 ��) @8�Z$���?!             J@       �       �                 @3�@H%u��?              I@       �       �                   @C@@�0�!��?             A@       �       �                 �|Y>@ܷ��?��?             =@       �       �                  sW@�X�<ݺ?             2@        �       �                 pf�@      �?              @       ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     $@        �       �                    A@"pc�
�?             &@       �       �                 �&B@����X�?             @        ������������������������       �                      @        �       �                   �?@���Q��?             @        ������������������������       �                     �?        �       �                   �@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �                     0@        ������������������������       �                      @        ������������������������       �                     "@        �       �                 �|�=@����?�?            �F@       ������������������������       �                    �A@        �       �                    ?@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                    (@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     �?��XI��?o            `f@       �       �                   �<@��H�}�?<             Y@        �       �                   �8@      �?             8@        �       �                    �?�q�q�?             "@       �       �                 ���Q@؇���X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?z�G�z�?             .@       ������������������������       �                     (@        ������������������������       �                     @        �       �                  �>@�w�"w��?/             S@        �       �                 �|�?@�P�*�?             ?@        �       �                 0C�<@      �?              @       ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ���=@
;&����?             7@       �       �                    �?D�n�3�?             3@        �       �                   @G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @L@��S���?
             .@       �       �                   �G@���|���?             &@       �       �                 ��:@և���X�?             @        ������������������������       �                      @        �       �                   �C@���Q��?             @        ������������������������       �                      @        �       �                   �F@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �G@:	��ʵ�?            �F@       �       �                   �@@$�q-�?             :@       ������������������������       �                     *@        �       �                    �?8�Z$���?             *@        �       �                   �A@�q�q�?             @        ������������������������       �                     �?        �       �                 @�Cq@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�����?             3@       �       �                    J@և���X�?
             ,@        �       �                 @�pX@؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    0@z\�3�?3            �S@        ������������������������       �                     @        �       �                     @DE��2{�?1            �R@        �       �                    �?������?             >@        ������������������������       �                     (@        �       �                    �?X�<ݚ�?	             2@        �       �                    *@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        �       �                    :@����X�?             @        ������������������������       �                     @        �       �                   P@@      �?             @        ������������������������       �                     �?        �       �                   �>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �                          �?:	��ʵ�?             �F@        �       �                    9@����X�?             5@        ������������������������       �                     @        �       �                 ��q1@և���X�?             ,@        ������������������������       �                     @        �       �                 03�7@���Q��?             $@        �       �                 �|�;@r�q��?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �T)D@      �?             @        ������������������������       �                     �?                               �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                              ���4@�8��8��?             8@                                 �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                 �?P���Q�?             4@        ������������������������       �                     @        	                      ���A@@4և���?             ,@        
                      ��T?@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������M}<���?g�/��?R0���[�?��)�?�3�=l}�?�\"<)H�?�q�q�?9��8���?              �?      �?        _�_�?���?�h
���?�~Y���?X`��?��~���?d!Y�B�?��7��M�?              �?      �?      �?              �?      �?                      �?�������?�������?      �?        �{a���?������?F]t�E�?/�袋.�?�������?�������?              �?UUUUUU�?�������?      �?      �?      �?      �?              �?      �?                      �?              �?      �?                      �?�?<<<<<<�?      �?                      �?�(\����?�G�z�?������?(������?{�G�z�?�z�G��?      �?      �?d!Y�B�?ӛ���7�?              �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?F]t�E�?]t�E�?      �?                      �?      �?              �?        �������?�?�q�q�?�q�q�?�؉�؉�?;�;��?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?9��8���?�q�q�?۶m۶m�?�$I�$I�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?      �?                      �?�?wwwwww�?۶m۶m�?I�$I�$�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?�.�袋�?F]t�E�?      �?        ��y��y�?�a�a�?      �?              �?      �?      �?      �?              �?      �?              �?        �*4��?��W�/��?�ҵ8f�?�iQR?δ?      �?        ]p�\p��?}�}��?      �?        z:�גC�?/,FBi�?�q�q�?�q�q�?              �?�s�9��?�c�1Ƹ?xxxxxx�?�?�������?�������?              �?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?         s�n_Y�?g\�5�?��RJ)��?�Zk��ֺ??�>��?l�l��?9��8���?�q�q�?۶m۶m�?�$I�$I�?      �?                      �?      �?      �?      �?                      �?      �?        7a~W��?�#{���?      �?      �?              �?      �?        �������?�?۶m۶m�?�$I�$I�?              �?      �?        q�����?;ڼOq��?;�;��?;�;��?)\���(�?���Q��?ZZZZZZ�?�������?��=���?a���{�?��8��8�?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        /�袋.�?F]t�E�?�m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?      �?              �?      �?              �?        �������?333333�?      �?                      �?      �?        ��I��I�?l�l��?      �?        �������?�������?              �?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���#��?���}��?{�G�z�?
ףp=
�?      �?      �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�������?�������?              �?      �?        ���k(�?��k(��?�RJ)���?�Zk����?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�Mozӛ�?Y�B��?l(�����?(������?      �?      �?              �?      �?        �?�������?F]t�E�?]t�E]�?�$I�$I�?۶m۶m�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?��O��O�?l�l��?�؉�؉�?;�;��?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?        Q^Cy��?^Cy�5�?�$I�$I�?۶m۶m�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?              �?        ��jq��?h *�3�?              �?,�Œ_,�?O贁N�?wwwwww�?�?      �?        r�q��?�q�q�?F]t�E�?t�E]t�?              �?      �?        �$I�$I�?�m۶m��?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��O��O�?l�l��?�m۶m��?�$I�$I�?      �?        �$I�$I�?۶m۶m�?      �?        �������?333333�?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?ffffff�?�������?      �?        n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ[س=hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������                           /@H���I�?�           8�@                                    @4���C�?'            �P@                                �-]@���N8�?             5@       ������������������������       �        	             3@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?���Q��?            �F@        	       
                 P��+@�	j*D�?             *@        ������������������������       �                     @                                   �?և���X�?             @                                 �-@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                   �?     ��?             @@        ������������������������       �                     �?                                @3�4@r֛w���?             ?@        ������������������������       �                     @                                   @ȵHPS!�?             :@                                   @�θ�?             *@        ������������������������       �                     @                                   @      �?             @                               ��T?@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@               Z                    �?dݿ�`�?�           (�@               M                    �?䖪@���?s            �g@              .                    �?b�L�4��?R            �`@                )                 `�@1@�:pΈ��?#             I@        !       "                     @�q�q�?             "@        ������������������������       �                      @        #       $                 �|�7@؇���X�?             @        ������������������������       �                      @        %       (                    �?z�G�z�?             @        &       '                 ��%@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        *       -                 03�=@��Y��]�?            �D@        +       ,                     �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     B@        /       :                     �?��s����?/             U@        0       9                   �H@>���Rp�?             =@       1       8                 �̾w@p�ݯ��?
             3@       2       3                    <@�t����?	             1@        ������������������������       �                     �?        4       7                    �?      �?             0@       5       6                    C@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        ;       >                   �6@�2����?            �K@        <       =                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       L                    �?ףp=
�?             I@       @       K                 �|�=@ i���t�?            �H@       A       B                   �<@�חF�P�?             ?@        ������������������������       �                     $@        C       D                     @���N8�?             5@        ������������������������       �                     �?        E       F                 �|Y=@      �?             4@        ������������������������       �                     �?        G       H                 ���@���y4F�?
             3@        ������������������������       �                      @        I       J                   @@���|���?             &@       ������������������������       ����Q��?             $@        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     �?        N       S                    �?|��?���?!             K@       O       P                     @ 7���B�?             ;@        ������������������������       �                     @        Q       R                   0:@�nkK�?             7@       ������������������������       �                     6@        ������������������������       �                     �?        T       Y                 X��E@�>����?             ;@       U       V                 ���@HP�s��?             9@        ������������������������       �                     @        W       X                 ��(@�KM�]�?
             3@       ������������������������       �؇���X�?             ,@        ������������������������       �                     @        ������������������������       �                      @        [       �                     @t�ۘ��?&           �|@        \       �                 `f�S@v�����?�             i@       ]       f                    �?�|����?t             f@        ^       c                   �K@h�����?&             L@       _       b                   �;@@3����?$             K@        `       a                    :@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     G@        d       e                   �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        g       |                 `ff:@      �?N             ^@       h       i                 �|Y=@��S�ۿ?0            �R@        ������������������������       �                     7@        j       k                     �?4��?�?!             J@        ������������������������       �                     @        l       o                 �|�=@�*/�8V�?            �G@        m       n                    @      �?             @       ������������������������       �                      @        ������������������������       �                      @        p       {                   �*@Du9iH��?            �E@       q       r                   �@@�����H�?             ;@        ������������������������       �                     &@        s       t                   @A@     ��?
             0@        ������������������������       �      �?             @        u       v                 `f�)@�8��8��?             (@        ������������������������       �                     @        w       x                   @D@z�G�z�?             @        ������������������������       �                      @        y       z                   �G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �        
             0@        }       �                     �?�<ݚ�?            �F@       ~       �                   �B@>��C��?            �E@              �                   �A@���Q��?             9@       �       �                   �>@�X����?             6@       �       �                 `fF<@b�2�tk�?             2@       �       �                   �K@�θ�?             *@       �       �                   @G@      �?             @       �       �                 �|�<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        ������������������������       �                      @        �       �                 ���a@�8��8��?             8@       ������������������������       �                     *@        �       �                    @"pc�
�?             &@       �       �                 `D�c@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        �       �                   @B@`�J�4��?�            p@       �       �                 �|�=@b�����?�            �k@       �       �                   �;@��8����?w             h@       �       �                 �T�I@6�`��V�?K             _@       �       �                   �@������?J            �^@        �       �                   �4@�(�Tw��?            �C@        �       �                    �?�KM�]�?             3@        ������������������������       �                      @        ������������������������       �        	             1@        �       �                   �5@�G�z��?             4@        �       �                 ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    7@X�Cc�?
             ,@        �       �                 ��@r�q��?             @        ������������������������       �                     @        �       �                 �?$@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?              @        �       �                   �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �Y�@���Q��?             @        �       �                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �:@H��?"�?3             U@       �       �                   �2@�C��2(�?0            @S@        �       �                    �?��s����?             5@        �       �                   �0@      �?             @        ������������������������       �                     �?        �       �                    �?���Q��?             @       �       �                 �y�+@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?��S�ۿ?
             .@       �       �                 pf� @�C��2(�?             &@        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�h����?"             L@        �       �                    �?�r����?             .@       �       �                   �9@�C��2(�?	             &@       ������������������������       �                     "@        �       �                 pf(@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���9@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��Y��]�?            �D@       �       �                   �4@ ���J��?            �C@        �       �                 @3�@���N8�?             5@        �       �                 �?�@r�q��?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     .@        ������������������������       �                     2@        ������������������������       �                      @        �       �                    �?և���X�?             @       �       �                 �� @���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��L@ =[y��?,             Q@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                 pf�@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        �       �                    �?�i�y�?'            �O@        �       �                 pf�3@�t����?	             1@        �       �                   �.@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     G@        �       �                 ��� @�z�G��?             >@       �       �                   @@@      �?             0@        �       �                   �@      �?              @        �       �                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �?�@r�q��?             @        ������������������������       �                     �?        �       �                   �?@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   @@@      �?	             ,@       �       �                   �>@����X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���/@����X�?             @        ������������������������       �                     @        �       �                   @A@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �                       @3�@��?^�k�?            �A@                               �?�@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     8@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������Q�Ȟ���?^-n����?'�l��&�?m��&�l�?�a�a�?��y��y�?              �?      �?      �?              �?      �?        333333�?�������?;�;��?vb'vb'�?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?���{��?�B!��?              �?��N��N�?�؉�؉�?ى�؉��?�؉�؉�?      �?              �?      �?333333�?�������?      �?                      �?              �?      �?        � V�b�?�S��;�?�
br1�?6�;���?v���?���-�?�Q����?��Q���?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ������?8��18�?�������?�������?      �?                      �?              �?z��y���?�a�a�?�i��F�?GX�i���?^Cy�5�?Cy�5��?�������?�������?              �?      �?      �?333333�?�������?      �?                      �?      �?                      �?      �?        ��7�}��?� O	��?�������?�������?              �?      �?        �������?�������?/�����?����X�?�Zk����?��RJ)��?      �?        �a�a�?��y��y�?      �?              �?      �?              �?6��P^C�?(������?      �?        ]t�E]�?F]t�E�?333333�?�������?      �?              �?              �?        	�%����?{	�%���?h/�����?	�%����?              �?d!Y�B�?�Mozӛ�?              �?      �?        �Kh/��?h/�����?q=
ףp�?{�G�z�?      �?        �k(���?(�����?۶m۶m�?�$I�$I�?      �?              �?        ����r�?ܸT��?q=
ףp�?��Q��?t�E]t�?]t�E�?�$I�$I�?�m۶m��?h/�����?���Kh�?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?      �?      �?�������?�?      �?        �N��N��?ى�؉��?      �?        r1����?m�w6�;�?      �?      �?      �?                      �?qG�w��?w�qGܱ?�q�q�?�q�q�?      �?              �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?        9��8���?�q�q�?$�;��?qG�w��?333333�?�������?�E]t��?]t�E]�?�8��8��?9��8���?ى�؉��?�؉�؉�?      �?      �?      �?      �?              �?      �?                      �?      �?        �������?�������?      �?                      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?F]t�E�?/�袋.�?�������?�������?      �?                      �?      �?        |�{�{��?����?G���w��?�B�I .�?�������?UUUUUU�?B!��?���{��?G:l��F�?�On���?�o��o��?� � �?�k(���?(�����?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?%I�$I��?�m۶m��?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �<��<��?1�0��?]t�E�?F]t�E�?z��y���?�a�a�?      �?      �?      �?        �������?333333�?      �?      �?              �?      �?                      �?�������?�?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?              �?        �$I�$I�?۶m۶m�?�������?�?]t�E�?F]t�E�?      �?              �?      �?              �?      �?              �?      �?              �?      �?        8��18�?������?��-��-�?�A�A�?��y��y�?�a�a�?�������?UUUUUU�?      �?              �?      �?      �?              �?              �?        ۶m۶m�?�$I�$I�?333333�?�������?      �?                      �?              �?              �?�������?�������?�������?�������?      �?              �?      �?      �?              �?      �?�������?AA�?<<<<<<�?�?9��8���?�q�q�?      �?                      �?      �?              �?        ffffff�?333333�?      �?      �?      �?      �?      �?      �?      �?                      �?�������?UUUUUU�?      �?        �������?�������?              �?      �?              �?              �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?_�_��?�A�A�?]t�E�?F]t�E�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJnխphG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM#hjh))��}�(h,h/h0M#��h2h3h4hph<�h=Kub������                       �U�R@<C�`��?�           8�@                                  @��y���?�           8�@                                    @������?             A@        ������������������������       �                     (@                                   �?���|���?             6@        ������������������������       �                     @                                @3�4@      �?             0@        ������������������������       �                     @        	       
                    @z�G�z�?	             $@        ������������������������       �                     @                                ��T?@���Q��?             @                                  @      �?             @        ������������������������       �                     �?                                03�9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?               c                    �?�K,���?{           (�@               &                     @f.i��n�?l            �f@                                  �*@�}�+r��?0             S@                                ��Y)@�S����?             3@                                 �F@@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?                                   <@���Q��?             @        ������������������������       �                     �?                                  �B@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                  @E@0�)AU��?$            �L@       ������������������������       �                    �F@                !                    �?�8��8��?             (@        ������������������������       �                      @        "       %                    :@ףp=
�?             $@        #       $                    5@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        '       L                    �?      �?<             Z@       (       7                  ��@b����?#            �O@        )       *                    �?�+$�jP�?             ;@        ������������������������       �                     @        +       2                 P�@�q�q�?             8@        ,       -                    �?      �?              @        ������������������������       �                      @        .       /                 ���@�q�q�?             @        ������������������������       �                     �?        0       1                 �|Y:@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        3       4                 ��@      �?             0@       ������������������������       �                     $@        5       6                 �&B@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        8       ?                  �#@)O���?             B@        9       :                   �1@�θ�?	             *@        ������������������������       �                     �?        ;       <                 `�X!@r�q��?             (@        ������������������������       �                     @        =       >                  SE"@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        @       G                    �?8����?             7@        A       F                 �|Y6@�q�q�?             @       B       C                 �&�)@�q�q�?             @        ������������������������       �                     �?        D       E                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        H       I                 03�0@@�0�!��?	             1@       ������������������������       �                      @        J       K                    �?�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        M       b                    @���� �?            �D@       N       O                   �0@     ��?             @@        ������������������������       �                      @        P       Y                 �|Y=@r�q��?             8@        Q       T                    �?z�G�z�?             $@        R       S                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        U       V                    �?      �?              @        ������������������������       �                     @        W       X                 ���9@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        Z       a                    �?d}h���?	             ,@        [       \                 �|�=@      �?             @        ������������������������       �                      @        ]       ^                 hV}1@      �?             @        ������������������������       �                      @        _       `                 `fV6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        d       �                     �?��!�?           {@        e       �                  �?@�ț��*�?5            �W@       f       m                    �?ڡR����?             �H@        g       h                 ���=@�q�q�?             @        ������������������������       �                     @        i       j                  Y>@�q�q�?             @        ������������������������       �                     �?        k       l                  �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        n       o                   �<@�K��&�?            �E@        ������������������������       �                     @        p                          @=@�99lMt�?            �C@       q       r                 ��$:@>���Rp�?             =@        ������������������������       �                     "@        s       t                 03k:@��Q��?             4@        ������������������������       �                     @        u       ~                 `f�;@������?
             1@       v       }                   �J@����X�?	             ,@       w       |                    H@և���X�?             @       x       y                 �|�?@���Q��?             @        ������������������������       �                     �?        z       {                   �C@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|Y=@�z�G��?             $@        ������������������������       �                      @        �       �                 X�lK@      �?              @       �       �                   �>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���}<S�?             G@        �       �                 �|Y:@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                    A@ >�֕�?            �A@        �       �                 �|Y>@      �?             0@       ������������������������       �                     "@        �       �                   @K@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@        �       �                 03�@�&�;���?�             u@        ������������������������       �                     ?@        �       �                     @�TM���?�            0s@        �       �                    �?���(-�?.            @R@        ������������������������       �                     @        �       �                    &@�����?(            �P@        �       �                    5@�KM�]�?
             3@        ������������������������       ����Q��?             @        ������������������������       �                     ,@        �       �                   �@@@��8��?             H@       ������������������������       �                     :@        �       �                   @A@���7�?             6@        �       �                   �3@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     2@        �       �                    �?�����8�?�            @m@        �       �                   �6@�%^�?            �E@        �       �                   �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03�-@>A�F<�?             C@       �       �                 ���@     ��?             @@        ������������������������       �                     $@        �       �                 �� @��2(&�?             6@       �       �                   @@�S����?
             3@       �       �                 �|=@8�Z$���?             *@        ������������������������       �                     @        �       �                 �|�=@z�G�z�?             $@       ������������������������       �      �?              @        ������������������������       �                      @        �       �                 �|Y=@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�;@�q�q�?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    '@p^�AL�?�            �g@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                 pff?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 0�H@0�#�.^�?            `g@       �       �                   �:@�h�ഭ�?{            �f@        �       �                 @3�@ ��ʻ��?,             Q@       ������������������������       �                     C@        �       �                    �?(;L]n�?             >@       �       �                 0S5 @���7�?             6@        �       �                   �1@�8��8��?             (@        ������������������������       �r�q��?             @        ������������������������       �                     @        ������������������������       �        	             $@        ������������������������       �                      @        �       �                   �;@Ԫ2��?O            �\@        ������������������������       �                      @        �       �                    �?      �?N             \@        �       �                   `3@      �?             @@       �       �                    �?��a�n`�?             ?@       �       �                 �|Y=@ �Cc}�?             <@        ������������������������       �                      @        �       �                 ��(@ ��WV�?             :@       �       �                 ���@�X�<ݺ?             2@        ������������������������       �                     @        �       �                 X��A@@4և���?	             ,@       ������������������������       ��8��8��?             (@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �C@      �?;             T@       �       �                 `f�'@؇���X�?3            �Q@       �       �                 ��) @д>��C�?(             M@       �       �                 @3�@�*/�8V�?!            �G@       �       �                   @C@     ��?             @@       �       �                 �|Y>@��� ��?             ?@       �       �                 �|Y=@�8��8��?             8@        ������������������������       �                      @        �       �                  sW@�C��2(�?             6@        �       �                 pf�@r�q��?             (@       ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �                     $@        �       �                 �&B@����X�?             @        ������������������������       �                      @        �       �                   �?@���Q��?             @        ������������������������       �                     �?        �       �                   �A@      �?             @       �       �                   �@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        �       �                 �|Y=@�eP*L��?             &@       �       �                 ���"@r�q��?             @        ������������������������       �                      @        �       �                   �<@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �̜!@z�G�z�?             @        ������������������������       �                      @        �       �                 �|�=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     $@                                  �?���Q��?             @                             �|�;@�q�q�?             @        ������������������������       �                     �?                              �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                 �?     ��?*             P@              	                   �?r٣����?            �@@       ������������������������       �                     .@        
                        �4@X�<ݚ�?	             2@        ������������������������       �                     @                                 �?և���X�?             ,@                              �	U@�q�q�?             "@                               �}S@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                              �Vs@r�q��?             @                             @�pX@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 !@�n`���?             ?@        ������������������������       �                      @                                 �?\-��p�?             =@       ������������������������       �                     6@                                 �G@և���X�?             @                               �D@      �?             @                             ��n^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        !      "                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0M#KK��h2h3h4hVh<�h=Kub�������������܍�W�?/�F�JP�?-�Q���?ɥ�\���?�?xxxxxx�?              �?F]t�E�?]t�E]�?              �?      �?      �?              �?�������?�������?      �?        333333�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�~jmr�?1�+%�?�>�>��?�`�`�?(�����?�5��P�?^Cy�5�?(������?�$I�$I�?n۶m۶�?              �?      �?        �������?333333�?      �?              �?      �?              �?      �?        p�}��?��Gp�?              �?UUUUUU�?UUUUUU�?              �?�������?�������?�������?�������?              �?      �?                      �?      �?      �?�eY�eY�?5M�4M��?B{	�%��?/�����?              �?�������?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?�������?333333�?              �?      �?              �?      �?              �?UUUUUU�?�������?      �?                      �?��8��8�?9��8���?ى�؉��?�؉�؉�?              �?�������?UUUUUU�?      �?        �m۶m��?�$I�$I�?              �?      �?        8��Moz�?d!Y�B�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        �������?ZZZZZZ�?              �?UUUUUU�?UUUUUU�?              �?      �?        jW�v%j�?,Q��+�?      �?      �?      �?        UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        I�$I�$�?۶m۶m�?      �?      �?              �?      �?      �?      �?              �?      �?              �?      �?              �?              �?        �E��ģ�?��V}�p�?�~�-q��?�a�+�?����S��?����X�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?��)kʚ�?���)k��?              �?5H�4H��?�o��o��?�i��F�?GX�i���?      �?        �������?ffffff�?              �?xxxxxx�?�?�m۶m��?�$I�$I�?۶m۶m�?�$I�$I�?333333�?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        333333�?ffffff�?      �?              �?      �?      �?      �?              �?      �?                      �?ӛ���7�?d!Y�B�?/�袋.�?F]t�E�?              �?      �?        ��+��+�?�A�A�?      �?      �?      �?        �m۶m��?�$I�$I�?      �?                      �?      �?        �9J���?3�E��?      �?        �j�Z�?���/�?��իW��?�P�B�
�?      �?        g��1��?���@��?�k(���?(�����?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?        �.�袋�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?        �������?���?�}A_��?�}A_�?�������?�������?      �?                      �?������?Cy�5��?      �?      �?      �?        ��.���?t�E]t�?(������?^Cy�5�?;�;��?;�;��?      �?        �������?�������?      �?      �?      �?        �������?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?i�O{�?��)_�%�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��b���?w��?-�-��?�~�~�?�������?�?      �?        �������?�?�.�袋�?F]t�E�?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?              �?              �?        $���>��?p�}��?              �?      �?      �?      �?      �?�s�9��?�c�1Ƹ?%I�$I��?۶m۶m�?              �?O��N���?;�;��?��8��8�?�q�q�?      �?        n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?              �?              �?                      �?      �?      �?۶m۶m�?�$I�$I�?a���{�?|a���?r1����?m�w6�;�?      �?      �?�{����?�B!��?UUUUUU�?UUUUUU�?      �?        ]t�E�?F]t�E�?�������?UUUUUU�?      �?        333333�?�������?      �?        �m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        t�E]t�?]t�E�?�������?UUUUUU�?      �?              �?      �?      �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?      �?|���?>���>�?              �?�q�q�?r�q��?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �c�1��?�9�s��?      �?        �{a���?a����?              �?�$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�[�.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K���h2h3h4hph<�h=Kub��������       N                 ���$@�,�٧��?�           8�@                                   �?���c���?�            @p@               
                    �?�p ��?            �D@                                ���@      �?             0@        ������������������������       �                     �?                                 s�@��S�ۿ?             .@        ������������������������       �                     @               	                    �?�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?                                 sW@�+e�X�?             9@                                ���@�q�q�?             @        ������������������������       �                     �?                                pf�@���Q��?             @                                �|Y:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 �#@�KM�]�?
             3@                               `�X!@�X�<ݺ?	             2@        ������������������������       �                     $@                                  �;@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?               K                    �?���;QU�?�            `k@                                   @P�p�(+�?�            �j@        ������������������������       �                      @               8                 �|Y=@����$�?�            �i@                5                   �<@���z�k�?A            �Y@       !       4                   �;@<����?<            �W@       "       %                    �?�5U��K�?5            �T@        #       $                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        &       +                 @3�@p`q�q��?3            �S@       '       *                 ���@�&=�w��?"            �J@        (       )                  Md@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     E@        ,       3                   �:@���B���?             :@       -       2                 pf� @      �?             8@        .       1                   �3@      �?             (@        /       0                   �1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             (@        ������������������������       �                      @        ������������������������       �                     (@        6       7                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        9       >                    �?��9J���?C             Z@        :       =                   @@�IєX�?	             1@       ;       <                 ���@�8��8��?             (@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ?       @                    �?�d���?:            �U@        ������������������������       �        
             1@        A       B                   �?@��?^�k�?0            �Q@        ������������������������       �                     @@        C       D                 �&B@�}�+r��?             C@        ������������������������       �                     0@        E       F                 P�@�C��2(�?             6@        ������������������������       �                     �?        G       J                 @3�@���N8�?             5@        H       I                   �A@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             0@        L       M                ��k!@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        O       z                    �?ڀ���?           0|@        P       [                    �?p�|����?H            @\@       Q       R                     @`Jj��?'             O@       ������������������������       �                     E@        S       Z                 `�@1@z�G�z�?             4@       T       W                    �?�	j*D�?             *@       U       V                 �|Y6@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        X       Y                 �|Y=@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        \       y                   @J@j���� �?!            �I@       ]       n                     �?�s��:��?             C@       ^       _                 ��2>@ �o_��?             9@        ������������������������       �                     @        `       g                 X�,@@�q�q�?             5@        a       f                 �|Y;@�eP*L��?             &@       b       e                   �8@r�q��?             @       c       d                 0wff@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        h       m                    C@ףp=
�?             $@        i       l                    �?z�G�z�?             @       j       k                   �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        o       t                   �5@�θ�?             *@        p       s                    �?�q�q�?             @       q       r                 �y.@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        u       v                 �|Y=@ףp=
�?	             $@       ������������������������       �                     @        w       x                     @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        {       �                    B@�F�*i��?�             u@       |       �                     @��?��?�            �n@       }       �                    �?     ��?Z             b@       ~                           �? ��N8�?1             U@        ������������������������       �                     �?        �       �                    �?��'�`�?0            �T@       �       �                   �;@@�E�x�?            �H@        �       �                   �:@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     C@        ������������������������       �                     A@        �       �                    �?������?)             N@       �       �                    :@�{��?��?&             K@        �       �                     �?�X�<ݺ?             2@        ������������������������       �                      @        �       �                    &@      �?             0@        �       �                    5@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �        
             *@        �       �                 ��yC@�E��ӭ�?             B@       �       �                   @A@J�8���?             =@       �       �                   �@@�n_Y�K�?             :@       �       �                     �?8����?             7@       �       �                   @>@և���X�?             ,@        �       �                 �|Y=@r�q��?             @        ������������������������       �                     @        �       �                 `f�;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|�<@      �?              @        ������������������������       �                     @        �       �                   �>@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 `fF)@�����H�?             "@        ������������������������       �                     @        �       �                 �|Y<@z�G�z�?             @        ������������������������       �                      @        �       �                 �|�=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    *@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���1@�کd�?@            �Y@        �       �                    �?���Q��?             D@       �       �                 ���.@� �	��?             9@        �       �                 �|�=@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                 �|�;@�q�q�?             .@        ������������������������       �                     @        �       �                    �?r�q��?	             (@       �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�r����?             .@       �       �                    �?؇���X�?             ,@       �       �                   �*@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��Y7@���N8�?(            �O@        �       �                    �?�ՙ/�?             5@       �       �                 �|�7@�q�q�?             (@       �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 03C3@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�����H�?             "@        �       �                 м�5@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��T?@r�q��?             E@       �       �                    �?���7�?             6@        �       �                 �|�:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        �       �                 ��p@@�z�G��?             4@        ������������������������       �                     @        �       �                 �T�I@��S�ۿ?
             .@        ������������������������       �                     "@        �       �                    �?r�q��?             @        �       �                    ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�����?;            �V@        ������������������������       �                      @        �       �                     �?ؤ�u��?7            �T@        �       �                    @@      �?             @@        �       �                    �?�q�q�?             "@        ������������������������       �                     @        �       �                 `fF<@      �?             @        �       �                    J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?\X��t�?             7@        ������������������������       �                     @        �       �                    J@�E��ӭ�?             2@       �       �                  x#J@�eP*L��?             &@        ������������������������       �                     @        �       �                 ���a@      �?              @       �       �                   �B@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��[�8��?!            �I@        �       �                     @ҳ�wY;�?             1@       �       �                    L@�θ�?	             *@       �       �                   @F@�C��2(�?             &@        �       �                   �E@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   @C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     A@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub��������������&��jq�?:�g *�?;�;��?�;�;�?dp>�c�?8��18�?      �?      �?      �?        �?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        R���Q�?���Q��?UUUUUU�?UUUUUU�?              �?�������?333333�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�k(���?(�����?��8��8�?�q�q�?      �?              �?      �?      �?                      �?              �?�ܹs���?�1bĈ�?��C���?^�
�u��?      �?        3y����?j6��bP�?���O ��?ch���V�?���%N�?�X�0Ҏ�?���h��?��k���?      �?      �?              �?      �?        T:�g *�?^-n����?tHM0���?�x+�R�?/�袋.�?F]t�E�?      �?                      �?      �?        ��؉���?ى�؉��?      �?      �?      �?      �?      �?      �?      �?                      �?      �?              �?                      �?      �?              �?      �?              �?      �?        ;�;��?�؉�؉�?�?�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        �:���C�?Ȥx�L��?      �?        _�_��?�A�A�?      �?        �5��P�?(�����?      �?        ]t�E�?F]t�E�?              �?��y��y�?�a�a�?�������?�������?      �?                      �?      �?              �?      �?              �?      �?        `����_�?P� 	P�?04��A�?h�e�&_�?�B!��?���{��?              �?�������?�������?;�;��?vb'vb'�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?                      �?�������?ZZZZZZ�?�k(���?��k(��?�Q����?
ףp=
�?              �?UUUUUU�?UUUUUU�?t�E]t�?]t�E�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?�������?�������?�������?      �?      �?              �?      �?                      �?              �?ى�؉��?�؉�؉�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?�������?�������?      �?              �?      �?      �?                      �?      �?        ���]�`�?	j*D>�?���/>�?u)���?      �?      �?�a�a�?�y��y��?              �?��k���?1P�M��?9/���?և���X�?F]t�E�?]t�E�?              �?      �?                      �?              �?wwwwww�?�?���^B{�?/�����?��8��8�?�q�q�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?              �?        �q�q�?r�q��?�rO#,��?|a���?;�;��?ى�؉��?d!Y�B�?8��Moz�?�$I�$I�?۶m۶m�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?333333�?�������?              �?      �?        �q�q�?�q�q�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        UUUUUU�?�������?              �?      �?        ��,��?��6��;�?�������?333333�?�Q����?)\���(�?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�?�������?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�a�a�?��y��y�?�<��<��?�a�a�?�������?�������?�������?�������?      �?                      �?�$I�$I�?۶m۶m�?      �?                      �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?        �������?UUUUUU�?�.�袋�?F]t�E�?      �?      �?      �?                      �?      �?        ffffff�?333333�?              �?�������?�?      �?        �������?UUUUUU�?      �?      �?              �?      �?              �?        h�h��?�/��/��?      �?        4u~�!��?�%���?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?              �?      �?                      �?!Y�B�?��Moz��?              �?�q�q�?r�q��?t�E]t�?]t�E�?      �?              �?      �?UUUUUU�?�������?      �?                      �?      �?              �?        �?�������?�������?�������?�؉�؉�?ى�؉��?F]t�E�?]t�E�?�������?�������?              �?      �?                      �?      �?              �?      �?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��=hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM#hjh))��}�(h,h/h0M#��h2h3h4hph<�h=Kub������       �                 pF�,@���*1�?�           8�@               i                 `f�$@.�mQ��?�            �t@                                  �?�w>�
��?�             o@               	                   �3@      �?             D@                                �&B@ףp=
�?             $@                               �?@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        
                        �̌@��S���?             >@                                  �?      �?             4@                                  �?r�q��?             2@                               ���@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@                                pff@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                @3�@ףp=
�?	             $@                                  �8@�q�q�?             @        ������������������������       �                     �?                                �?�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                    @�`�k�?�             j@        ������������������������       �                     $@               .                    �?P���+�?|            �h@               -                   @@     ��?             @@              &                   �6@������?             ;@                !                 ��y@      �?              @        ������������������������       �                      @        "       #                 ���@r�q��?             @        ������������������������       �                      @        $       %                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        '       (                 ���@�KM�]�?	             3@        ������������������������       �                     (@        )       *                 �|�:@����X�?             @        ������������������������       �                     �?        +       ,                 �|�=@�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     @        /       F                   �:@�S-�?l            �d@        0       E                   @8@���7�?,            �P@       1       4                 ���@�1�`jg�?$            �K@        2       3                 �&b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        5       D                   �4@ ��WV�?"             J@       6       7                   �1@`Jj��?             ?@        ������������������������       �                     $@        8       C                 0S5 @�����?             5@       9       >                   �2@8�Z$���?	             *@        :       =                    �?�q�q�?             @       ;       <                 ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ?       @                 �?�@ףp=
�?             $@        ������������������������       �                     @        A       B                 @3�@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     5@        ������������������������       �                     &@        G       `                 ��) @�_�s���?@            @Y@       H       I                 ���@����\�?:            �V@        ������������������������       �                     6@        J       O                    �?ДX��?-             Q@        K       N                 X�I@ףp=
�?
             4@       L       M                 ��(@�t����?	             1@       ������������������������       �      �?             0@        ������������������������       �                     �?        ������������������������       �                     @        P       U                 �|Y>@8��8���?#             H@       Q       R                 �|Y=@�g�y��?             ?@        ������������������������       �                     @        S       T                  sW@`2U0*��?             9@        ������������������������       �      �?             @        ������������������������       �                     5@        V       _                   �C@������?             1@       W       Z                   �@���Q��?	             $@        X       Y                 �&B@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        [       \                   �?@����X�?             @        ������������������������       �                     �?        ]       ^                   �B@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        a       b                 ��y @�eP*L��?             &@        ������������������������       �                     @        c       h                   �>@      �?              @       d       g                   �<@���Q��?             @       e       f                   �;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        j       �                     @ҳ�wY;�?5            @U@       k       l                    �?�&�5y�?(             O@        ������������������������       �                     �?        m       x                    �?�'N��?'            �N@        n       w                   �J@     ��?             0@       o       p                 ��Y)@�r����?             .@        ������������������������       �                      @        q       r                    :@����X�?             @        ������������������������       �                     �?        s       t                   �A@r�q��?             @       ������������������������       �                     @        u       v                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        y       �                 �|�=@�:�^���?            �F@        z       �                    �?"pc�
�?             6@       {       �                 �|�<@z�G�z�?             4@       |                           &@�����H�?             2@        }       ~                    5@      �?              @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     7@        �       �                 0S�*@\X��t�?             7@        ������������������������       �                     &@        �       �                    �?r�q��?             (@       �       �                   �4@      �?              @        �       �                   �-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �A@��T��?�            �w@       �       �                    �?2��8c�?�            �o@        �       �                   �>@ �&�T�?6             W@       �       �                    �?�G�z.�?0             T@        �       �                    �?��<D�m�?            �H@       �       �                    �?@4և���?             E@       ������������������������       �                     5@        �       �                     @؇���X�?	             5@        ������������������������       �                     @        �       �                    @d}h���?             ,@       �       �                  S�2@      �?              @       �       �                 �|Y=@���Q��?             @       �       �                    3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                  "&d@�g�y��?             ?@       �       �                 �|Y<@X�<ݚ�?             ;@        �       �                    �?����X�?             ,@       �       �                 pV�C@�C��2(�?             &@        ������������������������       �                     @        �       �                    8@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��.@�n_Y�K�?             *@        ������������������������       �                      @        �       �                 �|�=@���!pc�?	             &@       �       �                  �v6@�q�q�?             "@        ������������������������       �                     @        �       �                    �?���Q��?             @       �       �                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        �       �                 03SA@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �RL@      �?             (@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?
;&����?b             d@       �       �                    @�q�q�?4            @T@        ������������������������       �                     @        �       �                     @ �o_��?1            �R@       �       �                    �?��<b�ƥ?             G@        �       �                    <@P���Q�?             4@        �       �                     �?r�q��?             @        ������������������������       �                     @        �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                     :@        �       �                 ��Y1@8^s]e�?             =@        �       �                    9@      �?              @        ������������������������       �                     @        �       �                 �|�;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?؇���X�?             5@        ������������������������       �                      @        �       �                 `fV6@�S����?             3@        ������������������������       �                     �?        �       �                    @�����H�?             2@        ������������������������       �                      @        ������������������������       �        
             0@        �       �                    #@���Q8�?.             T@        �       �                   �C@�d�����?             3@       �       �                 @3�4@      �?	             0@       ������������������������       �                     $@        �       �                     @�q�q�?             @        ������������������������       �                     @        �       �                 @3;:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �9@f>�cQ�?#            �N@        ������������������������       �        
             2@        �       �                 `ff:@RB)��.�?            �E@        ������������������������       �        
             2@        �       �                    �?��H�}�?             9@       �       �                   �<@�û��|�?             7@        �       �                      @؇���X�?             @        ������������������������       �                     @        �       �                    ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|Y>@     ��?
             0@       ������������������������       �                     *@        ������������������������       �                     @        ������������������������       �                      @        �                           @��C�ח�?L             _@       �                           �?4��@���??             Y@       �       �                   �D@      �?5            �T@        �       �                   @C@      �?             0@       �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        �       �                 03�Q@z�G�z�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                          �?�{r٣��?'            �P@        �                         �I@�����?             5@       �                          �?z�G�z�?             $@       �                          �?����X�?             @        �                        ��A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@                                �R@�<ݚ�?            �F@                                @@&^�)b�?            �E@              
                  �K@�eP*L��?
             &@              	                ��:@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                �H@     ��?             @@                              x#J@r�q��?	             2@        ������������������������       �                     "@                                 �?�q�q�?             "@                               �G@      �?              @                             0�nL@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                      @                                 �?�q�q�?
             2@                                 �?      �?              @                                D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@              "                  @C@�8��8��?             8@               !                   �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             .@        �*       h�h))��}�(h,h/h0M#KK��h2h3h4hVh<�h=Kub������������`l����??'��d�?J�����?�>Q=h��?%����?��k���?      �?      �?�������?�������?      �?      �?              �?      �?                      �?�������?�?      �?      �?UUUUUU�?�������?F]t�E�?]t�E�?      �?                      �?�$I�$I�?�m۶m��?      �?                      �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?        ��|z�?7c,�?      �?        ���/M�?�Q7���?      �?      �?B{	�%��?{	�%���?      �?      �?      �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?�k(���?(�����?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?              �?        ���A#��?J���冸?�.�袋�?F]t�E�?A��)A�?�־a�?UUUUUU�?UUUUUU�?      �?                      �?O��N���?;�;��?���{��?�B!��?      �?        =��<���?�a�a�?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �������?�������?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?              �?              �?        ��g����?Q`ҩy�?.؂-؂�?�>�>�?      �?        �������?ZZZZZZ�?�������?�������?<<<<<<�?�?      �?      �?      �?              �?        �������?�������?��{���?�B!��?      �?        ���Q��?{�G�z�?      �?      �?      �?        xxxxxx�?�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?                      �?      �?        ]t�E�?t�E]t�?              �?      �?      �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?�������?:�s�9�?�1�c��?      �?        �����?ާ�d��?      �?      �?�?�������?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        }�'}�'�?l�l��?/�袋.�?F]t�E�?�������?�������?�q�q�?�q�q�?      �?      �?      �?      �?      �?              �?                      �?      �?              �?        ��Moz��?!Y�B�?              �?�������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        1x]o<�?�C|Q�a�?Ely(���?�I��6�?���,d�?��7��M�?ffffff�?ffffff�?և���X�?��S�r
�?�$I�$I�?n۶m۶�?              �?�$I�$I�?۶m۶m�?              �?۶m۶m�?I�$I�$�?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?              �?�B!��?��{���?�q�q�?r�q��?�$I�$I�?�m۶m��?F]t�E�?]t�E�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        ;�;��?ى�؉��?              �?F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?              �?              �?      �?      �?                      �?Y�B��?�Mozӛ�?UUUUUU�?UUUUUU�?      �?        �Q����?
ףp=
�?d!Y�B�?��7��M�?�������?ffffff�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?|a���?	�=����?      �?      �?              �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?        (������?^Cy�5�?              �?�q�q�?�q�q�?              �?      �?        �������?ffffff�?y�5���?Cy�5��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��!XG�?�u�y���?      �?        S֔5eM�?���)k��?      �?        {�G�z�?
ףp=
�?8��Moz�?��,d!�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?      �?        [k���Z�?J)��RJ�?�(\����?�G�z�?      �?      �?      �?      �?�q�q�?r�q��?              �?�������?�������?      �?              �?      �?              �?      �?                      �?��|��?|���?�a�a�?=��<���?�������?�������?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?9��8���?�q�q�?���/��?�}A_��?t�E]t�?]t�E�?UUUUUU�?�������?      �?                      �?      �?              �?      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?�������?UUUUUU�?              �?      �?                      �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?9��8���?�q�q�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��(hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                 03�I@n��"�)�?�           8�@              �                    �?���r�Q�?r           ��@              <                    �?p�����?-           �|@               1                    .@"��$�?E            �[@              
                 ��@4�B��?/            �R@                                ���@�C��2(�?             6@        ������������������������       �                     $@               	                    �?r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @                                   �?
j*D>�?"             J@                                    @      �?              @        ������������������������       �                      @                                  �-@r�q��?             @                                  �,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               (                   @B@d�
��?             F@                                   @���|���?            �@@                                `f�)@�8��8��?             (@        ������������������������       �                     @                                   ;@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @               '                  �#@�G��l��?             5@              "                   �9@b�2�tk�?             2@              !                 xF� @z�G�z�?             $@                                 �2@      �?             @        ������������������������       �                     �?                                   �7@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        #       $                    ;@      �?              @        ������������������������       �                     @        %       &                 �|Y>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        )       0                     @"pc�
�?             &@       *       +                    D@      �?              @        ������������������������       �                     @        ,       /                   �'@���Q��?             @       -       .                   �J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        2       7                    �?������?            �B@        3       6                     �?�q�q�?             "@       4       5                   �H@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        8       9                    �?h�����?             <@        ������������������������       �                     @        :       ;                   �2@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        =       �                   @S@T���D9�?�            �u@       >       Y                    �?
���?�            �u@        ?       L                 �|Y=@RB)��.�?            �E@        @       K                 ��d8@�eP*L��?             &@       A       B                     @�q�q�?             "@        ������������������������       �                     �?        C       D                 ��@      �?              @        ������������������������       �                     �?        E       F                 ��Y&@և���X�?             @        ������������������������       �                     �?        G       H                 �0@�q�q�?             @        ������������������������       �                     �?        I       J                   �2@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        M       R                   `A@      �?             @@       N       Q                   @@ �q�q�?             8@        O       P                 ���@�C��2(�?             &@       ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �        	             *@        S       X                   `E@      �?              @        T       U                   �B@      �?             @        ������������������������       �                      @        V       W                      @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        Z       �                   @>@�t����?�             s@       [       v                     @������?�            �q@        \       ]                    @��O���?7            @U@        ������������������������       �                     (@        ^       a                     �?L������?/            @R@        _       `                   �<@؇���X�?             ,@        ������������������������       �                      @        ������������������������       �                     (@        b       u                   �*@�j��b�?(            �M@       c       t                   �F@�S����?             C@       d       i                 `fF)@z�G�z�?             >@        e       h                    5@�����H�?             "@        f       g                   �2@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        j       k                 �|�<@���N8�?             5@        ������������������������       �                      @        l       m                 �|�=@�n_Y�K�?             *@        ������������������������       �                     �?        n       s                   �C@�q�q�?             (@       o       p                    @@�<ݚ�?             "@        ������������������������       �                     @        q       r                   �A@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     5@        w       �                 ��Y @ܴD��?�            @i@       x       �                   �4@0�й���?c            @b@        y       ~                   �3@��+7��?             7@       z       {                 �?�@�	j*D�?             *@       ������������������������       �                     @        |       }                   �1@�q�q�?             @        ������������������������       �      �?              @        ������������������������       �      �?             @               �                 P�@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                 @3�@������?T            �^@       �       �                   �>@\�t��Y�?F            �Y@       �       �                   �8@@4և���?1            �Q@        �       �                 ���@8�Z$���?             *@        �       �                 ���@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �<@�}�+r��?&            �L@        ������������������������       �                     1@        �       �                 ��(@��(\���?             D@       �       �                    �?�LQ�1	�?             7@       �       �                 ���@z�G�z�?
             .@        ������������������������       �                     @        �       �                 �|Y=@���!pc�?             &@        ������������������������       �                     �?        ������������������������       �z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                     1@        �       �                    �?�'�`d�?            �@@        ������������������������       �                      @        �       �                   @@@��a�n`�?             ?@        �       �                   �?@      �?             $@        �       �                 pff@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 P�@և���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        �       �                   @C@�����?             5@        ������������������������       �                     &@        �       �                    D@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     4@        �       �                    �?h�����?#             L@        �       �                   `3@؇���X�?             @       ������������������������       �                     @        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���!@@�E�x�?            �H@        �       �                   �:@���N8�?             5@        ������������������������       �                     &@        �       �                 @Q!@ףp=
�?             $@        ������������������������       �                     @        �       �                 �|Y<@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@        �       �                   �>@D�n�3�?             3@        ������������������������       �                     @        �       �                   �B@8�Z$���?	             *@        �       �                 �|�<@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     @��%��?E            �[@        �       �                    �?<���D�?            �@@       ������������������������       �                     8@        �       �                    *@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    @���L��?0            �S@        �       �                    �?����"�?             =@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             8@        �       �                    @�C��2(�?             &@        ������������������������       �                     @        �       �                 @3�2@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @��
ц��?             *@       �       �                    @�q�q�?             (@       �       �                 `f�:@      �?             $@        ������������������������       �                     @        �       �                    @r�q��?             @        ������������������������       �                     @        �       �                 ��T?@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @�D��?            �H@       �       �                 �A7@v�X��?             F@       �       �                    �?�q�����?             9@        �       �                 03�-@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                    )@���Q��?	             .@        �       �                 ���4@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���!pc�?             &@        �       �                    <@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        ������������������������       �                     @        �       �                    �?��~٩�?Q            `a@       �       �                 �|�=@�x�E~�?1            @V@        �       �                 �|Y=@@4և���?             <@       ������������������������       �                     4@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �N@        �       
                   �?� �	��?              I@       �                            @�P�*�?             ?@       �       �                    �?�5��?             ;@       �       �                 p"�X@�n_Y�K�?	             *@       �       �                  �}S@      �?              @       ������������������������       �                     @        �       �                 0�HU@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 p�w@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 `f�K@և���X�?             ,@        ������������������������       �                      @        �                        �|Y>@�q�q�?             (@        ������������������������       �                      @                                �D@z�G�z�?             $@        ������������������������       �                     @                              ���[@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @                                 ;@      �?             @        ������������������������       �                     �?              	                �|�>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                 �?���y4F�?             3@                                �?�z�G��?             $@                             @�ys@����X�?             @                                B@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                 6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������o怖�?�� 3���?�y��3m�?��*�%�?�r�^��?B���?Nq��$�?�~G����?L�Ϻ��?�Y7�"��?F]t�E�?]t�E�?              �?UUUUUU�?�������?              �?      �?        ;�;��?b'vb'v�?      �?      �?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?�.�袋�?�袋.��?F]t�E�?]t�E]�?UUUUUU�?UUUUUU�?              �?�q�q�?�q�q�?      �?                      �?1�0��?��y��y�?�8��8��?9��8���?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?      �?      �?                      �?              �?/�袋.�?F]t�E�?      �?      �?      �?        333333�?�������?      �?      �?              �?      �?                      �?      �?        к����?��g�`��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?�$I�$I�?�m۶m��?              �?d!Y�B�?�Mozӛ�?      �?                      �?���NV��?��Ħ��?0�甹��?A�`���?S֔5eM�?���)k��?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?                      �?              �?      �?      �?�������?UUUUUU�?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?              �?      �?      �?              �?      �?              �?        <<<<<<�?�?�|����?������?�������?�?      �?        �Ǐ?~�?����?۶m۶m�?�$I�$I�?              �?      �?        �N��?��/���?(������?^Cy�5�?�������?�������?�q�q�?�q�q�?�������?�������?      �?              �?      �?      �?        �a�a�?��y��y�?      �?        ;�;��?ى�؉��?              �?UUUUUU�?UUUUUU�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?        �(0���?z��~�X�?����?����Ǐ�?zӛ����?Y�B��?vb'vb'�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?      �?�������?�������?      �?                      �?�|����?������?P ���E�?��VCӽ?n۶m۶�?�$I�$I�?;�;��?;�;��?      �?      �?      �?                      �?      �?        �5��P�?(�����?      �?        �������?333333�?��Moz��?Y�B��?�������?�������?      �?        F]t�E�?t�E]t�?              �?�������?�������?      �?              �?        6�d�M6�?'�l��&�?      �?        �c�1��?�s�9��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?�������?�������?=��<���?�a�a�?      �?        �������?�������?              �?      �?              �?        �m۶m��?�$I�$I�?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        և���X�?9/���?��y��y�?�a�a�?      �?        �������?�������?      �?        �������?�������?              �?      �?              �?        l(�����?(������?              �?;�;��?;�;��?333333�?�������?              �?      �?              �?                      �?}���g�?���L�?|���?|���?              �?�q�q�?r�q��?              �?      �?        �4H�4H�?��o��o�?�i��F�?	�=����?�������?�������?              �?      �?        �������?�������?F]t�E�?]t�E�?              �?UUUUUU�?�������?              �?      �?        �؉�؉�?�;�;�?�������?�������?      �?      �?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ������??4և���?�.�袋�?颋.���?���Q��?�p=
ף�?333333�?ffffff�?      �?                      �?333333�?�������?      �?      �?              �?      �?        F]t�E�?t�E]t�?      �?      �?              �?      �?              �?              �?              �?        p�l�:��?��$D��?p�\��?����G�?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?                      �?�Q����?)\���(�?�Zk����?�RJ)���?/�����?h/�����?ى�؉��?;�;��?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?                      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?6��P^C�?(������?ffffff�?333333�?�m۶m��?�$I�$I�?�������?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���~hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM)hjh))��}�(h,h/h0M)��h2h3h4hph<�h=Kub������       �                     @� ��4d�?�           8�@               S                     �?���Ɉ��?�            �r@              $                    �?,Tg�x��?e             e@                                ��<J@     ��?*             P@                                   �?"pc�
�?             &@                                03�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        	       
                 �|�;@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @               #                    �?`��}3��?"            �J@                                 @E@�D��?             �H@                                  �?     ��?             @@       ������������������������       �                     6@                                   �?      �?             $@                                 �5@      �?              @        ������������������������       �                      @                                Ȫ�c@�q�q�?             @        ������������������������       �                     @                                X�,@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   >@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?��.k���?
             1@        ������������������������       �                     @                                м�M@z�G�z�?             $@        ������������������������       �                     �?               "                 �U�T@�����H�?             "@                !                 xCQ@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        %       J                   �J@z0��k��?;             Z@       &       -                    �?�0���?1            �T@        '       (                 ���a@ �#�Ѵ�?            �E@       ������������������������       �                    �@@        )       *                    �?z�G�z�?             $@        ������������������������       �                     @        +       ,                 Ъ�c@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        .       I                    �?�Q����?             D@       /       H                    �?��J�fj�?            �B@       0       =                   `@@��.k���?             A@        1       <                    F@����X�?	             ,@       2       ;                   @>@X�<ݚ�?             "@       3       4                 �̌*@և���X�?             @        ������������������������       �                     �?        5       :                 �|�?@      �?             @       6       7                 �|Y=@      �?             @        ������������������������       �                     �?        8       9                 `fF<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        >       ?                  x#J@�z�G��?             4@        ������������������������       �                     "@        @       A                 �|Y>@�eP*L��?             &@        ������������������������       �                     @        B       G                 ��9L@      �?              @       C       D                   �C@      �?             @        ������������������������       �                     �?        E       F                    G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        K       P                 `��R@؇���X�?
             5@       L       O                   �R@�����H�?             2@       M       N                    �?�IєX�?             1@        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     �?        Q       R                   �O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        T       �                  I?@��rq���?^            �`@       U       t                 �|�=@��\j���?U            �^@        V       q                    �?T����1�?*             M@       W       X                    �?D�n�3�?             C@        ������������������������       �                     @        Y       d                   �;@      �?             @@       Z       _                    &@p�ݯ��?             3@        [       \                    �?      �?              @        ������������������������       �                     @        ]       ^                    5@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        `       c                    �?"pc�
�?
             &@        a       b                   �7@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        e       f                 `f&'@�	j*D�?	             *@        ������������������������       �                      @        g       h                 `f�)@"pc�
�?             &@        ������������������������       �                     @        i       p                   �7@      �?              @       j       k                    �?�q�q�?             @        ������������������������       �                      @        l       o                    1@      �?             @       m       n                 �|�<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        r       s                   �(@R���Q�?             4@        ������������������������       �                     @        ������������������������       �                     1@        u       �                    @     ��?+             P@       v       �                    �?r֛w���?*             O@        w       �                    �?r�q��?             2@       x       �                   �7@     ��?             0@       y       �                   �*@�r����?             .@       z       {                    �?"pc�
�?             &@        ������������������������       �                     �?        |                          �'@z�G�z�?             $@        }       ~                   �J@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    B@r�q��?             @        ������������������������       �                     @        �       �                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @A@`���i��?             F@        �       �                    �?�}�+r��?             3@        ������������������������       �                     @        �       �                   �@@��S�ۿ?
             .@       ������������������������       �                     &@        �       �                   �3@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     9@        ������������������������       �                      @        �       �                    �?"pc�
�?	             &@       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?rC���e�?�            �y@        �       �                    �?�2�R�?F            @^@        �       �                    @ �o_��?             I@       �       �                    �?�D��?            �H@        �       �                 `�@1@���Q��?             .@       �       �                    (@�	j*D�?             *@        ������������������������       �                     @        �       �                 �%@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �0@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @;@H�V�e��?             A@        �       �                    '@�q�q�?             "@        ������������������������       �                     �?        �       �                    -@      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @       �       �                 83*@z�G�z�?             @       �       �                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �|�=@`2U0*��?             9@       �       �                 �|=@�IєX�?
             1@        ������������������������       �                     @        �       �                    �?@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?DX�\��?)            �Q@        �       �                    @\-��p�?             =@       ������������������������       �                     9@        ������������������������       �                     @        �       �                    �?�����?             E@       �       �                  ��@<���D�?            �@@        ������������������������       �                      @        �       �                 ��(@�J�4�?             9@       �       �                 �|Y=@"pc�
�?             6@        ������������������������       �                      @        �       �                 X�I@ףp=
�?             4@       ������������������������       ������H�?
             2@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �       �                 �?�@�N5X��?�            r@        �       �                    �?��<D�m�?=            �X@       �       �                 P�J@�*v��?<            @X@        ������������������������       �                     ;@        �       �                   �@�#-���?+            �Q@       �       �                   �4@(L���?            �E@        ������������������������       �                     $@        �       �                 P�N@"pc�
�?            �@@       �       �                    7@�����H�?             ;@        �       �                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|�<@�}�+r��?	             3@        ������������������������       �                     $@        �       �                 ��@�����H�?             "@        ������������������������       �                     @        �       �                 �|Y>@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    =@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ;@        ������������������������       �                     �?        �       �                    �?�P��Af�?w            �g@        �       �                    �?f.i��n�?            �F@        �       �                 Ь�#@      �?             $@        �       �                   �8@z�G�z�?             @        ������������������������       �                     @        �       �                 03�!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 03�1@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ���4@��R[s�?            �A@        �       �                   �:@      �?              @       ������������������������       �                     @        �       �                    >@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 ��p@@�����H�?             ;@       �       �                    �?�θ�?
             *@        ������������������������       �                     @        �       �                 ��T?@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        �                       @3�@b<g���?X            @b@        �                          :@�eP*L��?             &@        �                          �4@z�G�z�?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @                                �A@r�q��?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @                                 $@�r����?Q            �`@                              @3�4@X�<ݚ�?             2@        ������������������������       �                     @              	                   �?�C��2(�?             &@       ������������������������       �                      @        
                         @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @              (                   �?lZ�?��?E            @]@                                3@8��8���?9             X@                              ��Y @�	j*D�?             *@                                 1@�q�q�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @              #                �T)D@�+Ĺ+�?3            �T@             "                   ?@@-�_ .�?/            �R@                             ��) @HP�s��?"             I@        ������������������������       �                     0@                              pf� @�t����?             A@        ������������������������       �                     �?              !                `�X#@�C��2(�?            �@@                              �|�=@r�q��?             2@                               �:@      �?             0@       ������������������������       �                     "@                                �;@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             .@        ������������������������       �                     8@        $      %                   ;@�<ݚ�?             "@        ������������������������       �                     �?        &      '                �|�>@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        �*       h�h))��}�(h,h/h0M)KK��h2h3h4hVh<�h=Kub��������������`uv��?,J>��?'Z��}�?p��(��?b�a��?��<��<�?      �?      �?/�袋.�?F]t�E�?      �?      �?      �?                      �?�q�q�?�q�q�?              �?      �?        M0��>��?�琚`��??4և���?������?      �?      �?              �?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?�?�������?              �?�������?�������?              �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?              �?        �;�;�?'vb'vb�?"�%��?o4u~�!�?�}A_Ч?�/����?              �?�������?�������?              �?�$I�$I�?�m۶m��?      �?                      �?�������?ffffff�?�"�u�)�?к����?�������?�?�$I�$I�?�m۶m��?�q�q�?r�q��?�$I�$I�?۶m۶m�?      �?              �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?ffffff�?333333�?      �?        ]t�E�?t�E]t�?      �?              �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?۶m۶m�?�$I�$I�?�q�q�?�q�q�?�?�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ����?&���g��?�����?�d����?�rO#,��?�FX�i��?(������?l(�����?              �?      �?      �?^Cy�5�?Cy�5��?      �?      �?              �?      �?      �?      �?      �?      �?        /�袋.�?F]t�E�?      �?      �?      �?                      �?      �?        ;�;��?vb'vb'�?      �?        F]t�E�?/�袋.�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?333333�?333333�?      �?                      �?      �?      �?���{��?�B!��?UUUUUU�?�������?      �?      �?�?�������?F]t�E�?/�袋.�?              �?�������?�������?      �?      �?              �?      �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?      �?                      �?F]t�E�?F]t�E�?�5��P�?(�����?      �?        �������?�?      �?              �?      �?              �?      �?              �?                      �?F]t�E�?/�袋.�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?6)[��5�?)[��5)�?��ˠ�?a���i��?
ףp=
�?�Q����?������??4և���?333333�?�������?vb'vb'�?;�;��?      �?        r�q��?�q�q�?              �?      �?      �?              �?      �?                      �?iiiiii�?ZZZZZZ�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ���Q��?{�G�z�?�?�?      �?        n۶m۶�?�$I�$I�?      �?                      �?      �?                      �?�]�����?�D+l$�?�{a���?a����?              �?      �?        =��<���?�a�a�?|���?|���?      �?        �z�G��?{�G�z�?/�袋.�?F]t�E�?              �?�������?�������?�q�q�?�q�q�?      �?              �?              �?        ]�l� �?�"�O�|�?��S�r
�?և���X�?���AG�? tT����?      �?        �A�A�?_�_�?⎸#��?w�qG��?      �?        /�袋.�?F]t�E�?�q�q�?�q�q�?      �?      �?              �?      �?        �5��P�?(�����?      �?        �q�q�?�q�q�?      �?        �������?�������?      �?      �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?              �?        + �-��?T��Iw�?�`�`�?�>�>��?      �?      �?�������?�������?      �?              �?      �?              �?      �?        �������?�������?              �?      �?        X|�W|��?PuPu�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?ى�؉��?�؉�؉�?      �?        �$I�$I�?۶m۶m�?      �?                      �?      �?        ֫W�^��?�P�B�
�?]t�E�?t�E]t�?�������?�������?UUUUUU�?UUUUUU�?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?�������?�?r�q��?�q�q�?              �?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?        =�C=�C�?^�^�?�������?�������?vb'vb'�?;�;��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        (፦ί�?���ˊ��?S�n0E�?к����?q=
ףp�?{�G�z�?      �?        <<<<<<�?�?              �?]t�E�?F]t�E�?�������?UUUUUU�?      �?      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?                      �?      �?              �?        9��8���?�q�q�?              �?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJCLUhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �6       K��R�}�(hKhiK�hjh))��}�(h,h/h0K煔h2h3h4hph<�h=Kub��������       ^                     @�t����?�           8�@                                   �?�h��?�             t@                                  �E@�?�0�!�?T             a@                                  �?P����?E            �]@              
                 ��*@ �ׁsF�?;             Y@                                `f�)@P���Q�?             4@        ������������������������       �                      @               	                    :@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �        -             T@                                p"$X@�X�<ݺ?
             2@       ������������������������       �                     ,@                                   $@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?r�q��?             2@                                   �?d}h���?             ,@                               ��A@ףp=
�?             $@                                ���;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   5@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               Q                     �?6zg�K��?m            @g@              N                    �?f�Sc��?;            �X@              %                   �<@P�%f��?7            �V@                                   �4@���!pc�?             &@        ������������������������       �                      @        !       "                 `f�D@�����H�?             "@        ������������������������       �                     @        #       $                   �;@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        &       M                 p�w@�J�j�?0            �S@       '       L                   �R@���!pc�?/            @S@       (       K                   @J@��{�?6�?.            �R@       )       J                    �?V��z4�?$             O@       *       7                  Y>@^n����?"             N@        +       6                   `G@��
ц��?             :@       ,       -                 03:@���|���?             6@        ������������������������       �                     @        .       /                 �|Y=@��S���?             .@        ������������������������       �                     @        0       1                 `f&;@���!pc�?             &@       ������������������������       �                     @        2       3                    �?և���X�?             @        ������������������������       �                     �?        4       5                 X��B@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        8       =                  x#J@H�V�e��?             A@       9       <                    �?P���Q�?             4@        :       ;                    C@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        >       ?                 �|Y>@և���X�?	             ,@        ������������������������       �                      @        @       C                    �?      �?             (@        A       B                   �H@      �?             @        ������������������������       �                      @        ������������������������       �                      @        D       E                    A@      �?              @        ������������������������       �                      @        F       G                 `�iJ@�q�q�?             @        ������������������������       �                     �?        H       I                 03�U@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             *@        ������������������������       �                      @        ������������������������       �                      @        O       P                 �̰f@      �?              @       ������������������������       �                     @        ������������������������       �                     @        R       S                    #@��|���?2             V@        ������������������������       �                     $@        T       ]                   �*@ ��WV�?-            �S@       U       \                   �A@@4և���?             E@       V       [                   �@@H%u��?             9@       W       Z                    &@�nkK�?             7@       X       Y                   �5@��S�ۿ?
             .@        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     B@        _       �                 `f�%@��VI��?�            Px@       `       �                   �?@h��Q(�?�            �p@       a       z                    �?r֛w���?�             k@        b       q                 P��@\��_��?*            �Q@        c       p                    �?�J�4�?             9@       d       e                 ��y@�<ݚ�?             2@        ������������������������       �                      @        f       i                 ���@      �?             0@        g       h                 �|�9@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        j       o                    �?����X�?             @       k       l                   �5@�q�q�?             @        ������������������������       �                     �?        m       n                 �|�:@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     @        r       y                    �?nM`����?             G@       s       t                    �?�X���?             F@        ������������������������       �                     ;@        u       x                    �?�t����?             1@       v       w                 �|Y=@      �?             0@        ������������������������       �                     �?        ������������������������       �        
             .@        ������������������������       �                     �?        ������������������������       �                      @        {       �                    �?�@i����?X            @b@       |       �                    �?`����?W            �a@        }       ~                    3@
j*D>�?             :@        ������������������������       �                     @               �                 �|Y>@�X����?             6@       �       �                    ;@����X�?             5@       �       �                   �9@և���X�?
             ,@       �       �                 pff@���!pc�?             &@        �       �                 pf�@      �?             @        ������������������������       �                     �?        �       �                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�=@ 	��p�?E             ]@       �       �                    �?@-�_ .�?B            �[@       �       �                   �:@�1�`jg�?A            �[@       �       �                   �0@����e��?)            �P@        �       �                 pFD!@r�q��?             @        �       �                 pf�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        %             N@        �       �                 ��) @�Ra����?             F@       ������������������������       �                    �B@        �       �                 ��)"@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �>@���Q��?             @       �       �                 (Se!@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        "            �I@        �       �                    �?���6�?O            @^@        �       �                 03�:@">�֕�?            �A@       �       �                    �?��a�n`�?             ?@       �       �                   �,@�S����?             3@        ������������������������       �                     @        �       �                    �?�θ�?	             *@        �       �                 �0@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?ףp=
�?             $@       ������������������������       �                      @        �       �                   `3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 03�-@�q�q�?             (@        �       �                 P��+@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @       ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @2X��ʑ�?9            �U@        �       �                 `f�:@����X�?
             ,@       �       �                    @ףp=
�?             $@        �       �                 ��0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @        �       �                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?<ݚ�?/             R@       �       �                    5@�z�G��?             D@        ������������������������       �                     $@        �       �                    @���Q��?             >@       �       �                    �?      �?             8@       �       �                    �?X�<ݚ�?             2@       �       �                 ���*@�eP*L��?             &@        ������������������������       �                     �?        �       �                 ��Y.@      �?             $@        ������������������������       �                      @        �       �                 �|�;@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                 `fV6@և���X�?             @       �       �                   �;@z�G�z�?             @        ������������������������       �                      @        �       �                 `fv1@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 �|�:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?     ��?             @@       �       �                 �T)D@�<ݚ�?             2@       ������������������������       �        
             ,@        ������������������������       �                     @        �       �                    )@@4և���?
             ,@        ������������������������       �                     �?        ������������������������       �        	             *@        �)       h�h))��}�(h,h/h0K�KK��h2h3h4hVh<�h=Kub�������������G�+J>�?r%�k���?�.>9�?��h�`��?�����Ң?�������?'u_[�?�V'u�?{�G�z�?�G�z��?�������?ffffff�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?��8��8�?              �?      �?      �?      �?                      �?UUUUUU�?�������?۶m۶m�?I�$I�$�?�������?�������?      �?      �?              �?      �?                      �?      �?      �?              �?      �?                      �?�Gy��?�p�7��?����>�?������?�O��O��?�`�`�?t�E]t�?F]t�E�?      �?        �q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?        ^-n����?D�#{��?F]t�E�?t�E]t�?�K~���?7�i�6�?2�c�1�?�s�9��?�������?DDDDDD�?�;�;�?�؉�؉�?]t�E]�?F]t�E�?      �?        �������?�?      �?        t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?iiiiii�?ZZZZZZ�?ffffff�?�������?�q�q�?�q�q�?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?      �?      �?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?              �?                      �?              �?      �?      �?              �?      �?        F]t�E�?颋.���?              �?O��N���?;�;��?n۶m۶�?�$I�$I�?)\���(�?���Q��?�Mozӛ�?d!Y�B�?�������?�?              �?      �?              �?                      �?      �?              �?        ���k�2�?}�$(���?�Wc"=P�?z�rv��?���{��?�B!��?$Zas �?�K=��?�z�G��?{�G�z�?9��8���?�q�q�?      �?              �?      �?9��8���?�q�q�?              �?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?      �?              �?        zӛ����?C���,�?�E]t��?]t�E�?              �?<<<<<<�?�?      �?      �?              �?      �?                      �?      �?        X�^�z��?�B�
*�?�v�'��?$Zas �?b'vb'v�?;�;��?              �?�E]t��?]t�E]�?�m۶m��?�$I�$I�?�$I�$I�?۶m۶m�?F]t�E�?t�E]t�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?                      �?������?�{a���?S�n0E�?к����?A��)A�?�־a�?�>����?|���?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ]t�E]�?]t�E�?      �?        �$I�$I�?�m۶m��?              �?      �?              �?        333333�?�������?      �?      �?      �?                      �?      �?                      �?      �?        =;n,��?���#���?�A�A�?_�_��?�s�9��?�c�1��?^Cy�5�?(������?              �?�؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        }A_���?}A_��?�$I�$I�?�m۶m��?�������?�������?      �?      �?              �?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?        �q�q�?��8��8�?ffffff�?333333�?      �?        333333�?�������?      �?      �?�q�q�?r�q��?]t�E�?t�E]t�?              �?      �?      �?      �?              �?      �?      �?                      �?۶m۶m�?�$I�$I�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?9��8���?�q�q�?      �?                      �?n۶m۶�?�$I�$I�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       P                  �#@S*f���?�           8�@                                   �?6"�MB�?�            �p@                                 SE"@r�z-��?!            �J@                                  �?�������?             F@              
                    �?�����?             5@              	                 ���@P���Q�?             4@                                0��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     �?                                  �@8����?             7@                                ��@؇���X�?             ,@                               �|Y:@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                   4@X�<ݚ�?             "@        ������������������������       �                     �?                                  �9@      �?              @        ������������������������       �                     @                                �?�@���Q��?             @        ������������������������       �                     �?                                �|�;@      �?             @        ������������������������       �                      @                                �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@               O                    �?��g�?�            @k@              N                   �?@tCo���?�            �j@               !                     @�C��2(�?c            �d@        ������������������������       �                      @        "       -                    �?P��-�?^            �c@        #       ,                   @@8�Z$���?             :@       $       '                   �6@r�q��?             8@        %       &                 ��y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        (       )                 �|=@��2(&�?	             6@        ������������������������       �                      @        *       +                 ���@d}h���?             ,@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                      @        .       G                 ���"@�1����?Q            ``@       /       D                   �>@0{�v��?M            @_@       0       7                 �|Y=@hx<?v��?K            �]@       1       2                 @3�@ ��PUp�?0            �Q@       ������������������������       �        #            �J@        3       6                   �2@�X�<ݺ?             2@        4       5                 ��Y @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             ,@        8       A                 ��) @8��8���?             H@       9       @                 �|�=@���}<S�?             G@       :       ?                 �Y5@������?            �D@       ;       >                 ��@8�Z$���?             :@       <       =                 ���@P���Q�?             4@       ������������������������       �                     (@        ������������������������       �      �?              @        ������������������������       �      �?             @        ������������������������       �        	             .@        ������������������������       �                     @        B       C                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        E       F                 pff@      �?             @        ������������������������       �                     @        ������������������������       �                     @        H       M                 �|�=@�q�q�?             @       I       L                 �|Y=@z�G�z�?             @       J       K                   �6@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        "            �H@        ������������������������       �                     @        Q       �                 03[L@�d�f���?           �{@       R       �                    @f?8���?�            �u@       S       t                 �B,@�i#[��?�             u@        T       e                    �?�f7�z�?2            �U@       U       d                   �J@ףp=
�?             I@       V       a                    �?      �?             H@       W       X                 pF%@`Ӹ����?            �F@        ������������������������       �                     &@        Y       `                   �9@�IєX�?             A@        Z       [                 �&�%@      �?              @        ������������������������       �                     �?        \       ]                 ��y)@؇���X�?             @       ������������������������       �                     @        ^       _                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     :@        b       c                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        f       g                    )@�MI8d�?            �B@        ������������������������       �                     @        h       i                 �|Y=@�FVQ&�?            �@@        ������������������������       �                     *@        j       k                 `fF)@ףp=
�?             4@        ������������������������       �                      @        l       s                   �*@r�q��?             (@       m       n                 �|�=@      �?              @        ������������������������       �                     �?        o       p                    B@؇���X�?             @        ������������������������       �                     @        q       r                   �F@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        u       �                     @�����?�             o@       v       �                    �?��.w��?S            `a@       w       �                    �?z�):���?=             Y@        x       {                     �?ȵHPS!�?             :@        y       z                 hލC@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        |       �                   �E@�t����?             1@       }       �                   �;@@4և���?	             ,@        ~                          �9@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     �?|�U&k�?-            �R@       �       �                   �J@<|ۤ$�?!            �K@       �       �                   �B@�ݏ^���?            �F@       �       �                 �|�<@�!���?             A@        ������������������������       �                     @        �       �                    �?��>4և�?             <@        �       �                 ���<@���|���?             &@       �       �                 ��";@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �T!@@j���� �?             1@       �       �                   �G@����X�?
             ,@       �       �                 03:@X�<ݚ�?             "@        ������������������������       �                      @        �       �                 `fF<@����X�?             @       �       �                 X�,@@���Q��?             @        ������������������������       �                     �?        �       �                 03k:@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     $@        ������������������������       �                     3@        �       �                 ��Y=@:�&���?            �C@       �       �                   @A@���}<S�?             7@       ������������������������       �                     4@        �       �                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 �D C@     ��?             0@       �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                 ��@@r�q��?             @        ������������������������       �                      @        �       �                    0@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�X����?J            �[@        ������������������������       �                     @        �       �                    �?�e�}|�?H            �Z@        �       �                    �?��S���?"            �F@        �       �                 03�1@�����?             3@       �       �                    �?������?             1@        �       �                    �?؇���X�?             @        �       �                   �-@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �D@�z�G��?             $@       �       �                 @3�/@      �?              @        ������������������������       �                      @        �       �                   �0@r�q��?             @       �       �                 �|�;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 �A7@�	j*D�?             :@       �       �                 03�-@�q�q�?             (@        ������������������������       �                      @        �       �                   �0@�z�G��?	             $@       �       �                    �?���Q��?             @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @3�2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?@4և���?
             ,@        ������������������������       �                     @        �       �                    @�C��2(�?             &@        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?��.��?&            �N@       �       �                  �v6@(N:!���?            �A@       �       �                 ��d2@`2U0*��?             9@       ������������������������       �        
             1@        �       �                 ��`3@      �?              @        �       �                   �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03�7@�z�G��?             $@        ������������������������       �                     �?        �       �                 �T)D@�<ݚ�?             "@        ������������������������       �                     @        �       �                    ;@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�θ�?             :@       �       �                    �?���y4F�?             3@        ������������������������       �                     @        �       �                 032@      �?
             0@        �       �                 `ff/@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                 ��T?@����X�?             @        ������������������������       �                     @        �       �                 pf�C@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        �                           @�5��
J�?B             W@       �                         �L@�<ݚ�?@            �V@       �       �                    �?@�0�!��?<            @U@       �       �                    �? pƵHP�?"             J@       ������������������������       �                     E@        �       �                    $@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �                        03�M@4���C�?            �@@        ������������������������       �                     @                                 �?      �?             <@                                �?\X��t�?             7@                             p"�X@�eP*L��?             &@                             xCQ@�q�q�?             @        ������������������������       �                     �?                                �8@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        	      
                �̾w@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                �@@�q�q�?	             (@        ������������������������       �                     @                                 �?X�<ݚ�?             "@                                �?      �?              @        ������������������������       �                     �?                                �D@����X�?             @        ������������������������       �                     @                              ��#[@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?                                 6@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������H�7�?=�o�a��?�3���?��3����?�琚`��?����!�?/�袋.�?t�E]t�?�a�a�?=��<���?�������?ffffff�?      �?      �?              �?      �?                      �?      �?        8��Moz�?d!Y�B�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?r�q��?�q�q�?              �?      �?      �?      �?        �������?333333�?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        ���T��?���[��?
�N]���?�_���?]t�E�?F]t�E�?      �?        6��(S��?R��fu�?;�;��?;�;��?�������?UUUUUU�?      �?      �?      �?                      �?��.���?t�E]t�?      �?        I�$I�$�?۶m۶m�?      �?              �?      �?      �?        J�eDP�?����?V-��?;�O��n�?>�b>�b�?���Щ?��ۥ���?��V،?      �?        ��8��8�?�q�q�?      �?      �?              �?      �?              �?        �������?�������?ӛ���7�?d!Y�B�?�|����?������?;�;��?;�;��?ffffff�?�������?      �?              �?      �?      �?      �?      �?              �?              �?      �?              �?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?      �?                      �?      �?              �?        �k߰��?yJ���?p��f��? ��2)�?�a�a�?��<��<�?a���{�?O#,�4��?�������?�������?      �?      �?l�l��??�>��?              �?�?�?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        ��L���?L�Ϻ��?              �?>����?|���?      �?        �������?�������?      �?        �������?UUUUUU�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?        Cw�jXz�?z'*O�?!����?�:����?H�z�G�?q=
ףp�?�؉�؉�?��N��N�?�q�q�?�q�q�?      �?                      �?�?<<<<<<�?�$I�$I�?n۶m۶�?�������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�`�|��?E>�S��?��)A��?��7�}��?��I��I�?�[�[�?�������?�������?              �?I�$I�$�?۶m۶m�?F]t�E�?]t�E]�?�������?�������?              �?      �?                      �?ZZZZZZ�?�������?�$I�$I�?�m۶m��?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?�������?333333�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?              �?      �?              �?              �?              �?        �o��o��?�A�A�?d!Y�B�?ӛ���7�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?�E]t��?]t�E]�?              �?��V�9��?�R���?�?�������?^Cy�5�?Q^Cy��?�?xxxxxx�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?333333�?ffffff�?      �?      �?              �?UUUUUU�?�������?�������?�������?      �?                      �?              �?      �?              �?        vb'vb'�?;�;��?�������?�������?      �?        333333�?ffffff�?333333�?�������?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?n۶m۶�?�$I�$I�?      �?        ]t�E�?F]t�E�?      �?      �?      �?                      �?      �?        �����?������?|�W|�W�?�A�A�?���Q��?{�G�z�?      �?              �?      �?      �?      �?      �?                      �?      �?        ffffff�?333333�?              �?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?ى�؉��?�؉�؉�?6��P^C�?(������?              �?      �?      �?      �?      �?      �?                      �?      �?        �m۶m��?�$I�$I�?      �?              �?      �?              �?      �?              �?        �Mozӛ�?�,d!Y�?�q�q�?9��8���?�������?ZZZZZZ�?;�;��?'vb'vb�?              �?�������?�������?      �?                      �?'�l��&�?m��&�l�?              �?      �?      �?!Y�B�?��Moz��?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?                      �?�������?�������?      �?                      �?�������?�������?      �?        �q�q�?r�q��?      �?      �?      �?        �$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?      �?        �������?�������?              �?      �?              �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ"�a,hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       ^                    �?�����?�           8�@                                    �?���`��?�             i@                                   �?�!���?-             Q@                                 �H@�z�G��?!             I@                                  �?���@��?            �B@       ������������������������       �                     4@                                ���<@��.k���?             1@        ������������������������       �                     @        	       
                   �8@      �?	             (@        ������������������������       �                      @                                0�c@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?                                   J@��
ц��?	             *@        ������������������������       �                     @                                  �K@�q�q�?             "@        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                     @        ������������������������       �                     @                                hf$R@b�2�tk�?             2@                                  �:@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                  �e@�C��2(�?             &@        ������������������������       �                     @                                  �?@z�G�z�?             @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                /                 P��@�tL�|��?T            �`@        !       .                    �?�㙢�c�?             7@       "       -                    �?      �?             0@       #       $                 ��y@�q�q�?             (@        ������������������������       �                     �?        %       *                 ���@���|���?
             &@       &       '                    �?�q�q�?             "@        ������������������������       �                     �?        (       )                   �7@      �?              @        ������������������������       �                      @        ������������������������       �                     @        +       ,                 �|�8@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        0       G                    �?\�����?D            �[@       1       <                   �2@�2����?#            �K@        2       3                 P��+@����X�?             5@        ������������������������       �                     $@        4       9                    �?�eP*L��?             &@        5       8                 83C6@      �?             @       6       7                   �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        :       ;                    @և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        =       B                    �?l��\��?             A@        >       ?                 �|�<@�<ݚ�?             "@       ������������������������       �                     @        @       A                  S�2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        C       D                     @`2U0*��?             9@        ������������������������       �                      @        E       F                    �?�nkK�?             7@       ������������������������       �                     6@        ������������������������       �                     �?        H       S                 �|Y=@�rF���?!            �K@        I       L                    �?      �?	             0@        J       K                   �;@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        M       N                 �n6@�q�q�?             "@        ������������������������       �                      @        O       R                    �?؇���X�?             @        P       Q                    *@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       ]                 �|Y>@��-�=��?            �C@       U       \                    �?�J�4�?             9@       V       W                     @���}<S�?             7@        ������������������������       �                     @        X       Y                    �?ףp=
�?             4@        ������������������������       �                     @        Z       [                 ��(@�t����?             1@       ������������������������       �8�Z$���?             *@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@        _       �                    �?<q��F�?M           �@        `       y                     @�����?i            �c@       a       x                    �?���Lͩ�?5            �R@       b       c                     �?fP*L��?             F@        ������������������������       �                     1@        d       w                   �J@������?             ;@       e       p                   �B@z�G�z�?             9@       f       o                   �7@�����H�?             2@       g       l                    1@r�q��?	             (@       h       k                    :@ףp=
�?             $@        i       j                   �4@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        m       n                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        q       r                   �'@և���X�?             @        ������������������������       �                     @        s       v                    E@      �?             @       t       u                   �,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     ?@        z       �                    @F~��7�?4            �T@       {       �                    �?�o;����?1            �S@       |       �                 03�1@|��?���?$             K@       }       �                 `f�%@X�<ݚ�?            �F@       ~                          �3@X�Cc�?             <@        ������������������������       �                     @        �       �                    A@��<b���?             7@       �       �                 �|Y>@���N8�?             5@       �       �                 P�@z�G�z�?             4@        �       �                 �&B@�q�q�?             @       �       �                 ���@���Q��?             @       �       �                 pff@      �?             @       �       �                 �|Y:@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �*@�t����?             1@        ������������������������       �                     @        �       �                 �|�<@"pc�
�?             &@        �       �                    .@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �                 �|Y>@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @��H�}�?             9@        �       �                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �0@�d�����?
             3@        ������������������������       �                      @        �       �                 �|�:@�eP*L��?             &@       �       �                 ���9@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �                       0wkS@fP*L���?�             v@       �       �                     @�UQ��?�            �u@        �       �                    %@�)l�o��?N            @^@        ������������������������       �                     &@        �       �                 ��D:@X�;�^o�?I            �[@       �       �                   �*@���#�İ?)            �M@       �       �                    4@`Ӹ����?            �F@        �       �                    &@؇���X�?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        �       �                     �?P�Lt�<�?             C@        ������������������������       �                     @        �       �                    �?��?^�k�?            �A@       �       �                   �@@г�wY;�?             A@       ������������������������       �                     9@        �       �                   @A@�����H�?             "@        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                   �>@������?             �I@        �       �                   @C@
j*D>�?             :@        �       �                 �|Y=@r�q��?             @        �       �                 `fF<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `G@�z�G��?             4@        �       �                   �F@�����H�?             "@       �       �                   �E@r�q��?             @        ������������������������       �                     �?        ������������������������       �z�G�z�?             @        ������������������������       �                     @        �       �                    K@�eP*L��?             &@        ������������������������       �                     @        �       �                 `fF<@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �B@`2U0*��?             9@        �       �                   �A@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �       �                    #@hdpZ�L�?�            @l@        �       �                    @      �?             $@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @z�G�z�?             @       �       �                 (C45@�q�q�?             @        ������������������������       �                     �?        �       �                 ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �                          �?�`5���?�             k@       �                       �T)D@�P�U`��?~            `h@       �       �                 �?�@���8��?z            `g@        �       �                 ���@X;��?6            @V@        �       �                 �|�:@@�0�!��?             1@        �       �                  Md@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        +             R@        �       �                 0SE @�q��/��?D            �X@        �       �                   �3@�5��
J�?"             G@        �       �                    1@����X�?             @        ������������������������       �      �?              @        �       �                   �2@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        �       �                   �>@8�Z$���?            �C@       �       �                   �4@�����H�?             ;@        �       �                 @3�@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                 �|Y=@���}<S�?             7@        ������������������������       �                      @        �       �                 ��) @�r����?             .@       ������������������������       �        
             *@        ������������������������       �                      @        �       �                 @3�@      �?	             (@        �       �                   �?@և���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        ������������������������       �                     @        �                         �;@ pƵHP�?"             J@        �                       @�!@ ��WV�?             :@                                 � @�8��8��?             (@        ������������������������       �                     �?                                 8@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �        
             ,@        ������������������������       �                     :@                                 ;@      �?              @        ������������������������       �                     @        	      
                �|�>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�����������������?��܍��?�1����?*g��1�?�������?�������?333333�?ffffff�?к����?L�Ϻ��?              �?�?�������?      �?              �?      �?      �?        �������?�������?              �?      �?        �;�;�?�؉�؉�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        9��8���?�8��8��?۶m۶m�?�$I�$I�?              �?      �?        F]t�E�?]t�E�?              �?�������?�������?      �?      �?              �?      �?                      �?SKE,�?Z�iu���?�7��Mo�?d!Y�B�?      �?      �?UUUUUU�?UUUUUU�?      �?        ]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?              �?      �?              �?              �?        A��)A�?߰�k��?� O	��?��7�}��?�$I�$I�?�m۶m��?              �?t�E]t�?]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?۶m۶m�?              �?      �?        �������?------�?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?{�G�z�?���Q��?              �?d!Y�B�?�Mozӛ�?              �?      �?        yJ���?�־a��?      �?      �?�$I�$I�?�m۶m��?      �?                      �?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        }˷|˷�?�A�A�?�z�G��?{�G�z�?ӛ���7�?d!Y�B�?      �?        �������?�������?      �?        <<<<<<�?�?;�;��?;�;��?      �?                      �?      �?        &&&&&&�?�������?���JG�?�	�Z��?�K~��?�6�i�?]t�E]�?颋.���?              �?{	�%���?B{	�%��?�������?�������?�q�q�?�q�q�?UUUUUU�?�������?�������?�������?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?      �?      �?                      �?      �?              �?                      �?���ˊ��?��h���?�#{���?��	�Z�?{	�%���?	�%����?�q�q�?r�q��?%I�$I��?�m۶m��?              �?��,d!�?��Moz��?�a�a�?��y��y�?�������?�������?UUUUUU�?UUUUUU�?�������?333333�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?                      �?      �?        �?<<<<<<�?              �?F]t�E�?/�袋.�?      �?      �?              �?      �?                      �?�q�q�?�q�q�?      �?              �?      �?      �?                      �?{�G�z�?
ףp=
�?UUUUUU�?UUUUUU�?      �?                      �?Cy�5��?y�5���?      �?        t�E]t�?]t�E�?�$I�$I�?�m۶m��?              �?      �?              �?              �?        ]t�E�?��.���?�ba4{�?�wz.�?���!pc�?�T�x?r�?              �?�־a��?J��yJ�?��N��?'u_[�??�>��?l�l��?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        ���k(�?(�����?      �?        _�_��?�A�A�?�?�?      �?        �q�q�?�q�q�?      �?      �?      �?              �?              �?        xxxxxx�?�?b'vb'v�?;�;��?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?ffffff�?333333�?�q�q�?�q�q�?�������?UUUUUU�?      �?        �������?�������?      �?        t�E]t�?]t�E�?              �?۶m۶m�?�$I�$I�?      �?                      �?���Q��?{�G�z�?�������?�������?      �?                      �?      �?        ٠ɗ��?4��A�/�?      �?      �?�������?�������?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?��Kh/�?Lh/����?�����?����?o�W@�n�?�C�刴?�u�{���?�E(B�?ZZZZZZ�?�������?�$I�$I�?۶m۶m�?      �?                      �?      �?              �?        /����?և���X�?�,d!Y�?�Mozӛ�?�$I�$I�?�m۶m��?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?;�;��?;�;��?�q�q�?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?        ӛ���7�?d!Y�B�?      �?        �������?�?      �?                      �?      �?      �?�$I�$I�?۶m۶m�?              �?�������?�������?      �?        'vb'vb�?;�;��?O��N���?;�;��?UUUUUU�?UUUUUU�?      �?        ]t�E�?F]t�E�?      �?                      �?      �?              �?              �?      �?              �?�������?�������?      �?                      �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�8�hhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM!hjh))��}�(h,h/h0M!��h2h3h4hph<�h=Kub������       x                     @��t���?�           8�@               U                  x#J@����>��?�            ps@                                  @T�$@��?�            �j@        ������������������������       �                      @                                  �6@������?�            �i@                                   �?�����?            �H@       ������������������������       �                     9@                                   �?�q�q�?             8@       	       
                   �2@�q�q�?             .@       ������������������������       �                     @                                  �'@      �?             $@       ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �                     "@               R                   �@@��Y���?f            �c@              Q                   �?@̏�xQ��?U            �_@              P                    @��C�ח�?T             _@              I                   �K@|;�p)�?S            @^@                                  �?V�r��?I            @[@                                   �?�z�G��?
             $@                               `��,@�q�q�?	             "@        ������������������������       �                     �?                                  @@@      �?              @                                  �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?               ,                    �?4���C�??            �X@               %                   �2@������?            �B@              $                   �*@ �q�q�?             8@               !                   �B@�X�<ݺ?
             2@       ������������������������       �                     ,@        "       #                    D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        &       '                  �v7@�θ�?	             *@        ������������������������       �                     �?        (       )                    D@r�q��?             (@       ������������������������       �                     @        *       +                     �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        -       >                 ��D:@���-T��?)             O@       .       =                    1@Hm_!'1�?            �H@       /       0                 �|Y=@�J�4�?             9@        ������������������������       �                     "@        1       2                 �|�=@      �?             0@        ������������������������       �                     �?        3       4                 `fF)@z�G�z�?             .@        ������������������������       �                     @        5       <                   �F@�z�G��?             $@       6       ;                   �C@      �?              @       7       8                    @@z�G�z�?             @        ������������������������       �                     �?        9       :                   �A@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     8@        ?       @                    <@�n_Y�K�?
             *@        ������������������������       �                      @        A       H                   `H@���!pc�?	             &@       B       G                    �?z�G�z�?             $@       C       F                 `f�:@�<ݚ�?             "@        D       E                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        J       O                     �?�8��8��?
             (@        K       L                 `fF<@r�q��?             @       ������������������������       �                     @        M       N                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        S       T                    �?�חF�P�?             ?@        ������������������������       �                     @        ������������������������       �                     :@        V       g                 ���X@�q�Q�?=             X@       W       ^                    �?ףp=
�?&             N@       X       ]                     �?���N8�?             E@       Y       \                 0�"K@��Y��]�?            �D@        Z       [                 `�iJ@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �C@        ������������������������       �                     �?        _       `                    �?�<ݚ�?             2@       ������������������������       �                     (@        a       d                    �?�q�q�?             @        b       c                 03/O@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        e       f                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        h       s                    �?*O���?             B@       i       p                    �?      �?             6@       j       m                 X�,@@      �?
             0@        k       l                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        n       o                 ��)[@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        q       r                 �\@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        t       u                    �?؇���X�?
             ,@       ������������������������       �                     $@        v       w                 03c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        y       �                    �?�+e�X�?�             y@        z       �                 `v�6@Ć��H��?D            �Z@       {       �                    �?Ї?��f�?5            @U@        |       �                    �?      �?             D@        }       �                 �|Y=@և���X�?             5@       ~                          �0@�C��2(�?             &@       ������������������������       �                     @        �       �                 03�-@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?z�G�z�?             $@       �       �                    �?����X�?             @       �       �                 ��%@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y8@�}�+r��?             3@        ������������������������       �                     @        �       �                 ���@$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?�ݏ^���?            �F@       �       �                 ��&@�>$�*��?            �D@       �       �                   �3@�q�q�?             ;@        �       �                 �&B@      �?             @        �       �                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 @3�@��+7��?             7@       �       �                    ;@�eP*L��?             &@       �       �                   �9@؇���X�?             @        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        �       �                 03�1@X�Cc�?
             ,@       �       �                 ���*@      �?             (@        ������������������������       �                     @        �       �                 ��Y.@      �?              @        ������������������������       �                      @        �       �                 �|�;@r�q��?             @        �       �                    .@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��T?@���7�?             6@       ������������������������       �        	             &@        �       �                 ��p@@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    @�׺W4�?�            Pr@        �       �                    @X�<ݚ�?             "@       �       �                 �y�-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 �?�@`����?�            �q@        �       �                    �?     ��?S             `@        �       �                 �|Y=@r�q��?             2@        �       �                 ���@և���X�?             @        ������������������������       �                     @        �       �                   @8@      �?             @        ������������������������       �                      @        �       �                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             &@        �       �                    �?�1�`jg�?E            �[@       �       �                  ��@�X�<ݺ?D             [@        ������������������������       �                     F@        �       �                   �<@     ��?+             P@        ������������������������       �                     ;@        �       �                   �@�MI8d�?            �B@       �       �                 �|Y=@d}h���?             <@        ������������������������       �                     �?        �       �                    �?�+$�jP�?             ;@       �       �                 X��A@      �?             0@       ������������������������       ���S�ۿ?
             .@        ������������������������       �                     �?        �       �                   @@@���|���?             &@       �       �                 �&B@      �?              @       �       �                 �|Y>@�q�q�?             @       ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        �                         @@@Tݭg_�?_            �c@       �                          �?��ׂ�?P            ``@       �       �                    �?Ft����?I            �^@        �       �                    /@�z�G��?             $@        ������������������������       �                     @        �       �                    7@և���X�?             @        ������������������������       �                     �?        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �                       �|�=@d}h���?C             \@       �       �                 @�!@�\m����?<             Y@        �       �                   �3@^����?            �E@        �       �                   �1@��
ц��?             *@        �       �                   �0@      �?              @       ������������������������       �      �?             @        ������������������������       �                      @        �       �                 0S5 @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 ��) @r�q��?             >@       ������������������������       �                     4@        �       �                   �:@      �?             $@        ������������������������       �                     @        �       �                 �|Y<@r�q��?             @        ������������������������       �                     @        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                         �<@���5��?"            �L@       �       �                    �?@-�_ .�?            �B@       �       �                    9@`2U0*��?             9@       ������������������������       �        
             0@        �       �                    ;@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�8��8��?             (@        ������������������������       �                     @        �                        `f2@      �?              @        ������������������������       �                     �?        ������������������������       �                     @                                 �?      �?             4@                                `3@�q�q�?             @        ������������������������       �                      @                              03�7@      �?             @        ������������������������       �                      @        ������������������������       �                      @                              �|Y=@d}h���?             ,@        	      
                ���"@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@                                �?@�q�q�?             (@                                �>@z�G�z�?             @                             �̌!@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                              d�6@@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                 #@�����H�?             "@                              `f�9@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 �?`2U0*��?             9@        ������������������������       �                      @                                �B@�nkK�?             7@        ������������������������       �                     "@                               @3�@@4և���?             ,@        ������������������������       ��q�q�?             @        ������������������������       �                     &@        �*       h�h))��}�(h,h/h0M!KK��h2h3h4hVh<�h=Kub�������������nԾ���?5"W��6�?��f�?t�����?�b?-��?X:Ɂ���?      �?        ?���(�?ہ�v`��?����X�?^N��)x�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?�$I�$I�?�m۶m��?      �?                      �?�Ȟ��t�?-n����?�\.����?�F��h4�?[k���Z�?J)��RJ�?y?r����?�ˠT�?�,�M���?���d	l�?ffffff�?333333�?UUUUUU�?UUUUUU�?              �?      �?      �?۶m۶m�?�$I�$I�?              �?      �?                      �?      �?        m��&�l�?'�l��&�?к����?��g�`��?UUUUUU�?�������?�q�q�?��8��8�?              �?      �?      �?      �?                      �?              �?�؉�؉�?ى�؉��?      �?        UUUUUU�?�������?              �?�������?333333�?              �?      �?        [k���Z�?�RJ)���?Y�Cc�?9/���?�z�G��?{�G�z�?      �?              �?      �?              �?�������?�������?      �?        ffffff�?333333�?      �?      �?�������?�������?      �?              �?      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?              �?        ;�;��?ى�؉��?              �?F]t�E�?t�E]t�?�������?�������?9��8���?�q�q�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?                      �?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?              �?�Zk����?��RJ)��?              �?      �?        UUUUUU�?�������?�������?�������?�a�a�?��y��y�?������?8��18�?      �?      �?              �?      �?                      �?      �?        �q�q�?9��8���?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?      �?      �?      �?      �?�������?�������?              �?      �?        F]t�E�?/�袋.�?      �?                      �?�������?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        R���Q�?���Q��?!V��G&�?�S�rp��?�������?�������?      �?      �?۶m۶m�?�$I�$I�?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?�������?�������?�m۶m��?�$I�$I�?�������?UUUUUU�?              �?      �?                      �?      �?        (�����?�5��P�?              �?;�;��?�؉�؉�?      �?                      �?�[�[�?��I��I�?�18���?�����?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?                      �?zӛ����?Y�B��?]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?              �?        �m۶m��?%I�$I��?      �?      �?              �?      �?      �?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?                      �?�.�袋�?F]t�E�?      �?        ]t�E�?F]t�E�?              �?      �?        :f���M�?gB����?�q�q�?r�q��?UUUUUU�?UUUUUU�?              �?      �?                      �?�v�'��?$Zas �?     ��?      �?�������?UUUUUU�?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        A��)A�?�־a�?��8��8�?�q�q�?      �?              �?      �?      �?        ��L���?L�Ϻ��?I�$I�$�?۶m۶m�?              �?/�����?B{	�%��?      �?      �?�������?�?      �?        ]t�E]�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        � � �?�|˷|��?w�_�	)�?#����[�?�S\2��?C��6�S�?ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?                      �?I�$I�$�?۶m۶m�?�Q����?R���Q�?�qG��?w�qG��?�؉�؉�?�;�;�?      �?      �?      �?      �?      �?        �������?�������?              �?      �?        �������?UUUUUU�?      �?              �?      �?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?        �}��?��Gp�?S�n0E�?к����?���Q��?{�G�z�?      �?        �q�q�?�q�q�?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        I�$I�$�?۶m۶m�?      �?      �?      �?                      �?      �?        �������?�������?�������?�������?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?                      �?�q�q�?�q�q�?      �?      �?              �?      �?              �?        ���Q��?{�G�z�?      �?        �Mozӛ�?d!Y�B�?      �?        n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJP�dhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       D                     �?ʡ�;S��?�           8�@                                   �?o��Ա�?r            `i@                                   �? qP��B�?4            �U@                                  �?�}��L�?.            �R@                                03�=@h�����?             <@        ������������������������       �                     �?        ������������������������       �                     ;@        ������������������������       �                    �G@        	                        Ъ�c@�C��2(�?             &@        
                        ���[@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               '                    �?.��$�?>            @]@               "                   @H@
j*D>�?             J@                                  �?f���M�?             ?@                               ���<@      �?             8@        ������������������������       �                     @                                �|Y<@����X�?             5@        ������������������������       �                      @                                   C@��
ц��?             *@                               ��2>@���Q��?             $@        ������������������������       �                      @                                X�,@@      �?              @        ������������������������       �                     @                                @�Cq@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               !                   �?@����X�?             @                                  �4@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        #       &                   �H@�����?             5@        $       %                   �T@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     .@        (       A                    �?؇>���?%            @P@       )       :                   �B@��f/w�?#            �N@       *       9                    R@     ��?             @@       +       4                   �=@      �?             <@       ,       3                   �F@��2(&�?             6@       -       .                 03:@�z�G��?             $@        ������������������������       �                     @        /       0                 03k:@���Q��?             @        ������������������������       �                     �?        1       2                 X��B@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     (@        5       6                   �>@�q�q�?             @        ������������������������       �                     @        7       8                 �|�<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ;       <                    �? 	��p�?             =@        ������������������������       �                     �?        =       >                 03�T@@4և���?             <@       ������������������������       �                     9@        ?       @                  �6f@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        B       C                    @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        E       �                    �?l��э�?G           �@        F       �                    �?��P��?f            �d@       G       �                 м�9@fȮ�Б�?N            �_@       H       U                    �?X�Emq�?B            �Z@        I       R                    �?��P���?            �D@        J       M                    �?��
ц��?	             *@       K       L                   P,@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        N       O                 P��+@      �?             @        ������������������������       �                      @        P       Q                 83�0@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        S       T                 ���@@4և���?             <@        ������������������������       �                      @        ������������������������       �                     :@        V       {                   �?@^��>�b�?*            @P@       W       ^                     @"Ae���?             �G@        X       Y                   �'@����X�?             @        ������������������������       �                     @        Z       ]                    �?      �?             @       [       \                   �<@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        _       `                    @��Q���?             D@        ������������������������       �                     @        a       z                    �?���@��?            �B@       b       g                   �3@r֛w���?             ?@        c       f                   �2@      �?             @       d       e                 ��K)@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        h       q                 P�@z�G�z�?             9@        i       j                 pff@���Q��?             @        ������������������������       �                     �?        k       l                 ���@      �?             @        ������������������������       �                     �?        m       n                   �7@�q�q�?             @        ������������������������       �                     �?        o       p                 �&B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        r       w                 ��*@ףp=
�?
             4@       s       t                   �9@�X�<ݺ?             2@       ������������������������       �                     .@        u       v                 �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        x       y                 �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        |       }                   @B@�q�q�?
             2@        ������������������������       �                     @        ~       �                     @�eP*L��?             &@              �                   �,@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     5@        �       �                     @����>�?            �B@        ������������������������       �                     @        �       �                    �?ףp=
�?             >@        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��T?@@4և���?             <@       ������������������������       �        	             1@        �       �                 ��p@@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?�O�t]E�?�            �u@       �       �                     @H�����?�            �r@        �       �                 �|�=@�IєX�?-             Q@        �       �                    �?ףp=
�?             >@        ������������������������       �                     �?        �       �                    @ܷ��?��?             =@        ������������������������       �                     @        �       �                 �|Y=@��2(&�?             6@       �       �                    &@P���Q�?             4@        �       �                    8@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                      @        �       �                   �*@P�Lt�<�?             C@       �       �                   @D@�nkK�?             7@       ������������������������       �        	             .@        �       �                   �'@      �?              @        ������������������������       �                      @        �       �                   �F@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        	             .@        �       �                    ,@�h*����?�            �l@        ������������������������       �                     �?        �       �                   @@@�`"���?�            �l@       �       �                   �?@�חF�P�?y            @g@       �       �                   �:@��2(&�?r             f@        �       �                 ��q1@"pc�
�?7             V@       �       �                    �?��1��?4            �T@        �       �                 H�%@և���X�?             @       �       �                   �6@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 0S5 @���Lͩ�?0            �R@       �       �                 @3�@L紂P�?!            �I@       �       �                    �?���}<S�?             G@        ������������������������       �                     �?        �       �                 ���@�:�^���?            �F@        �       �                    7@      �?              @       ������������������������       �                     @        �       �                 �&b@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �4@@-�_ .�?            �B@        �       �                 �?�@"pc�
�?             &@       ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     :@        �       �                   �2@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     8@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                 �T)D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �<@�C��2(�?;             V@        ������������������������       �                     $@        �       �                 �|Y=@��-�=��?3            �S@        �       �                 �̌!@�q�q�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�=@�8��8��?/             R@       �       �                    �?�C��2(�?*            �P@        �       �                    �?`Jj��?             ?@        �       �                 p&�@ףp=
�?             $@       �       �                 ���@؇���X�?             @        ������������������������       �                      @        ������������������������       �z�G�z�?             @        ������������������������       �                     @        �       �                   `3@���N8�?             5@       ������������������������       �                     3@        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                  sW@(N:!���?            �A@        �       �                 pf�@�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �      �?             @        �       �                 ��) @$�q-�?             :@       ������������������������       �                     1@        �       �                 �̜&@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 d�6@@���Q��?             $@       �       �                   �@�q�q�?             @        ������������������������       �                     �?        �       �                 �?�@z�G�z�?             @        ������������������������       �                     �?        �       �                 ��I @      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?�@`���i��?             F@       ������������������������       �                     :@        �       �                 @3�@�X�<ݺ?             2@        ������������������������       ��q�q�?             @        ������������������������       �        	             .@        �                          �?���X�K�?!            �F@       �       �                     @��}*_��?             ;@        �       �                    6@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             8@        �       �                 ��}@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                  @�d�����?             3@                              03�6@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @                              032@$�q-�?	             *@                                �5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        	                         #@r�q��?             2@        
                         �?և���X�?             @        ������������������������       �                     �?                              pf�C@�q�q�?             @                                @�q�q�?             @        ������������������������       �                     �?                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������N���I5�?d�~`l��?��Gu��?"\E;�?�}A_З?��}A�?O贁N�?�_,�Œ�?�$I�$I�?�m۶m��?      �?                      �?              �?F]t�E�?]t�E�?�������?�������?              �?      �?                      �?�Y��Y��?�LɔL��?b'vb'v�?;�;��?��Zk���?��RJ)��?      �?      �?      �?        �$I�$I�?�m۶m��?              �?�؉�؉�?�;�;�?333333�?�������?              �?      �?      �?      �?              �?      �?      �?                      �?              �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?=��<���?�a�a�?UUUUUU�?UUUUUU�?              �?      �?              �?        �����? �����?XG��).�?��!XG�?      �?      �?      �?      �?��.���?t�E]t�?ffffff�?333333�?      �?        �������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?������?�{a���?      �?        n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        ��r�\.�?i4�F��?}���|�?������?��r�\.�?�F��h�?�}�	��?5�x+��?�����?������?�;�;�?�؉�؉�?�$I�$I�?۶m۶m�?              �?      �?              �?      �?              �?      �?      �?      �?                      �?�$I�$I�?n۶m۶�?      �?                      �?r#7r#7�?�����?�w6�;�?W�+���?�$I�$I�?�m۶m��?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?333333�?�������?              �?L�Ϻ��?к����?���{��?�B!��?      �?      �?333333�?�������?              �?      �?                      �?�������?�������?�������?333333�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?�������?��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?t�E]t�?]t�E�?�$I�$I�?�m۶m��?      �?                      �?      �?                      �?�u�)�Y�?���L�?              �?�������?�������?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?      �?        /�袋.�?F]t�E�?              �?      �?        �w�q�?��#�;�?�&��%�?��6@�Ҿ?�?�?�������?�������?      �?        ��=���?a���{�?      �?        ��.���?t�E]t�?ffffff�?�������?      �?      �?      �?      �?      �?              �?                      �?���k(�?(�����?�Mozӛ�?d!Y�B�?      �?              �?      �?      �?        �������?UUUUUU�?      �?      �?      �?              �?        �D�o-��?)�F@J��?              �?���aܯ�?m5x�@�?�Zk����?��RJ)��?��.���?t�E]t�?/�袋.�?F]t�E�?�+Q���?,Q��+�?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?        �6�i�?�K~��?�������?�������?ӛ���7�?d!Y�B�?      �?        }�'}�'�?l�l��?      �?      �?      �?              �?      �?      �?                      �?S�n0E�?к����?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?        �������?333333�?              �?      �?              �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?]t�E�?F]t�E�?      �?        }˷|˷�?�A�A�?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?]t�E�?F]t�E�?���{��?�B!��?�������?�������?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?        ��y��y�?�a�a�?      �?              �?      �?              �?      �?        |�W|�W�?�A�A�?9��8���?�q�q�?      �?              �?      �?�؉�؉�?;�;��?      �?        9��8���?�q�q�?              �?      �?              �?        �������?333333�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?F]t�E�?      �?        ��8��8�?�q�q�?UUUUUU�?UUUUUU�?      �?        l�l��?�'}�'}�?_B{	�%�?B{	�%��?UUUUUU�?UUUUUU�?              �?      �?              �?      �?�������?�������?      �?                      �?Cy�5��?y�5���?UUUUUU�?UUUUUU�?              �?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?UUUUUU�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�g?BhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM=hjh))��}�(h,h/h0M=��h2h3h4hph<�h=Kub������       �                     @S*f���?�           8�@               '                 ��/@�k���)�?�            �t@                                   @��|�	��?;            �V@        ������������������������       �                     "@               &                    �?���ȫ�?5            �T@              %                   �-@H���I�?3            �S@              $                 �J+@؀�:M�?0            �R@                                  &@��W3�?-            �Q@        	                           �?� �	��?             9@        
                          �J@�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @                                  �5@�8��8��?
             (@        ������������������������       �      �?              @        ������������������������       �                     $@                                �|Y<@8����?             G@        ������������������������       �                     .@               #                   @G@`՟�G��?             ?@                                 �(@���|���?             6@        ������������������������       �                     �?                                   �?�q�q�?             5@        ������������������������       �                     @                                   �?j���� �?             1@                                 �*@ףp=
�?             $@                                 �B@      �?              @       ������������������������       �                     @                                   D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                    @@؇���X�?             @        ������������������������       �                     @        !       "                   @B@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        (       �                   �K@�M�
FD�?�            `n@       )       ~                    �?"wO�a��?�            @k@       *       k                     �?:{hWXS�?y            �g@       +       T                 03/O@���j��?W            @a@       ,       7                    �?4�.�A�?,            �O@        -       .                 �|�;@�E��ӭ�?             2@        ������������������������       �                     @        /       6                    �?�q�q�?             .@       0       5                 �|�=@r�q��?
             (@        1       2                 �ܵ<@�q�q�?             @        ������������������������       �                     �?        3       4                 03SA@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        8       9                    7@��S���?            �F@        ������������������������       �                     @        :       ;                    �?և���X�?             E@        ������������������������       �                     $@        <       M                 �T!@@     ��?             @@       =       >                   �<@�q�q�?             .@        ������������������������       �                     @        ?       L                   @>@�eP*L��?
             &@       @       A                 ��:@      �?              @        ������������������������       �                     �?        B       G                 `f�;@և���X�?             @       C       D                 X��B@      �?             @        ������������������������       �                     �?        E       F                   @G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        H       I                 �|Y=@�q�q�?             @        ������������������������       �                     �?        J       K                 X��B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        N       O                   �;@������?
             1@        ������������������������       �                      @        P       Q                 0�J@�r����?	             .@       ������������������������       �                     &@        R       S                 �K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        U       \                   �8@�7�QJW�?+            �R@        V       W                    �?�n_Y�K�?             *@        ������������������������       �                     @        X       [                   �7@r�q��?             @        Y       Z                   �4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ]       ^                    �?��� ��?#             O@       ������������������������       �                     E@        _       d                 ��>Y@���Q��?             4@        `       a                    �?      �?              @       ������������������������       �                     @        b       c                   �D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        e       j                 p�w@�q�q�?             (@       f       g                    �?      �?              @        ������������������������       �                     @        h       i                 ���a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        l       m                    4@䯦s#�?"            �J@        ������������������������       �        
             *@        n       o                    �?      �?             D@        ������������������������       �                      @        p       y                    �?�\��N��?             C@       q       r                   �6@���>4��?             <@        ������������������������       �                     @        s       x                    �?\X��t�?             7@       t       u                   �E@@4և���?             ,@       ������������������������       �                     $@        v       w                   �H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        z       {                    <@�z�G��?             $@        ������������������������       �                     @        |       }                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @               �                    �?�>����?             ;@        �       �                    7@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     2@        �       �                    �?�+e�X�?             9@        �       �                    �?���Q��?             @       �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?R���Q�?
             4@       �       �                   @O@�θ�?             *@       �       �                   �M@�C��2(�?             &@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �                          �?X��"C�?�            �w@       �       �                 Ь�#@L� P?)�?�            0r@       �       �                 ��@�����?�            `n@        �       �                 ���@�~�4_��?<             V@       �       �                    �?X�;�^o�?(            �K@        �       �                    �?r�q��?             @       �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?@9G��?#            �H@        �       �                 ���@�C��2(�?             6@       �       �                   �7@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     &@        ������������������������       �                     ;@        �       �                 ��@���|���?            �@@        ������������������������       �                     �?        �       �                  ��@     ��?             @@        �       �                 �|Y;@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �|Y=@X�Cc�?             <@        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��s����?             5@       �       �                 X��A@���y4F�?             3@       �       �                    �?�	j*D�?	             *@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?M�D���?c            `c@        �       �                   �9@��
ц��?
             *@        ������������������������       �                     @        �       �                    ;@�q�q�?             "@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                 ��� @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �3@���J�?Y            �a@        �       �                   �1@�GN�z�?             6@        ������������������������       �                     @        �       �                   �2@�q�q�?             .@        �       �                 ��Y @����X�?             @       �       �                 ��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �?�@      �?              @        ������������������������       �                     @        �       �                 0S5 @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �:@��S�ۿ?N             ^@        �       �                   �4@�(\����?             D@        �       �                 @3�@�8��8��?             (@        �       �                 P�@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     <@        �       �                    �?p=
ףp�?7             T@        ������������������������       �                     @        �       �                   �;@���Lͩ�?2            �R@        �       �                 �� @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �<@����Q8�?0            �Q@        ������������������������       �                     $@        �       �                 �|Y=@��GEI_�?+            �N@        �       �                   `!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                  sW@����˵�?)            �M@        �       �                 �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��) @���U�?'            �L@       �       �                   �B@����?�?            �F@       ������������������������       �                    �B@        �       �                   �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�>@�8��8��?             (@        �       �                 �̜!@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                 ��Y)@�q�q��?"             H@        ������������������������       �                     @        �       �                    �?�L�lRT�?             �F@        �       �                    �?     ��?             0@        ������������������������       �                     @        �       �                 �|�;@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        �                          ;@ܷ��?��?             =@        �                           �?z�G�z�?             $@        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        �       �                 �0@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              �T)D@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                              �|�>@�}�+r��?             3@       ������������������������       �                     $@                              �T)D@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        	                         @t���D�?:            �U@        
                         �?X�Cc�?             <@        ������������������������       �                     @                                 @�q�q�?             8@                             @3�4@�G�z��?             4@        ������������������������       �                      @                              ���A@      �?             (@                                �?�q�q�?             "@        ������������������������       �                     @                                 @      �?             @        ������������������������       �                      @                              `f�:@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 �?      �?             @                                @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @              <                  @C@�BbΊ�?'             M@             5                `v�6@~���L0�?#            �H@             4                   @@���>4��?             <@              )                03�-@�q�����?             9@        !      "                ��!@z�G�z�?             $@        ������������������������       �                     @        #      $                  �#@�q�q�?             @        ������������������������       �                     �?        %      &                   �?z�G�z�?             @        ������������������������       �                     �?        '      (                  �;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        *      /                   �?������?             .@        +      .                   �?؇���X�?             @        ,      -                ���1@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        0      1                   7@      �?              @        ������������������������       �                     @        2      3                   �?���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        6      7                   �?�����?             5@        ������������������������       �                     �?        8      9                ��T?@ףp=
�?             4@        ������������������������       �                     "@        :      ;                X��@@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     "@        �*       h�h))��}�(h,h/h0M=KK��h2h3h4hVh<�h=Kub�������������H�7�?=�o�a��?��;���?�b@:��?�Q�Q�?�\��\��?      �?        �cp>��?28��1�?Q�Ȟ���?^-n����?E>�S��?v�)�Y7�?p�z2~��? �
���?�Q����?)\���(�?�؉�؉�?ى�؉��?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        d!Y�B�?8��Moz�?      �?        �1�c��?�s�9��?F]t�E�?]t�E]�?      �?        UUUUUU�?UUUUUU�?              �?ZZZZZZ�?�������?�������?�������?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?                      �?      �?                      �?;����?�s��w�?�߅���?�p=��?�"����?��2�|�?!Y�B�?ozӛ���?��i��i�?�,˲,��?r�q��?�q�q�?              �?UUUUUU�?UUUUUU�?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        �������?�?      �?        ۶m۶m�?�$I�$I�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?]t�E�?t�E]t�?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?xxxxxx�?�?              �?�������?�?      �?              �?      �?              �?      �?        0��b�/�?t�@�t�?ى�؉��?;�;��?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        �B!��?�{����?              �?�������?333333�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?      �?        �������?�������?              �?      �?                      �?�V�9�&�?�����?              �?      �?      �?      �?        �5��P�?y�5���?I�$I�$�?n۶m۶�?      �?        ��Moz��?!Y�B�?�$I�$I�?n۶m۶�?              �?      �?      �?      �?                      �?      �?        333333�?ffffff�?              �?333333�?�������?              �?      �?        h/�����?�Kh/��?�q�q�?9��8���?              �?      �?                      �?R���Q�?���Q��?�������?333333�?      �?      �?              �?      �?              �?        333333�?333333�?ى�؉��?�؉�؉�?]t�E�?F]t�E�?      �?      �?              �?      �?              �?                      �?      �?        �J�Y\�?\8�v���?Z�D�a��?���fy�?w�M���?�#*�6�?]t�E�?��.���?�־a��?J��yJ�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?������?9/���?]t�E�?F]t�E�?/�袋.�?F]t�E�?              �?      �?              �?              �?        ]t�E]�?F]t�E�?              �?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        %I�$I��?�m۶m��?�$I�$I�?۶m۶m�?              �?      �?        z��y���?�a�a�?6��P^C�?(������?vb'vb'�?;�;��?              �?      �?              �?              �?        =���?a�qa�?�;�;�?�؉�؉�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?      �?      �?                      �?A�6�?��RO�o�?�袋.��?]t�E�?      �?        UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?              �?      �?              �?      �?        �������?�?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?              �?        333333�?ffffff�?      �?        �6�i�?�K~��?      �?      �?      �?                      �?O�o�z2�?��Vج?      �?        �d����?;ڼOqɰ?      �?      �?      �?                      �?W'u_�?��/���?      �?      �?              �?      �?        	�#����?p�}��?��I��I�?l�l��?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?�I��I��?l�l��?      �?      �?              �?333333�?ffffff�?      �?                      �?��=���?a���{�?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?�5��P�?(�����?      �?        �q�q�?�q�q�?      �?                      �?�;⎸�?$�;��?�m۶m��?%I�$I��?              �?�������?�������?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?      �?              �?      �?              �?              �?      �?      �?      �?              �?      �?                      �?�{a��?���=��?����>4�?������?I�$I�$�?n۶m۶�?���Q��?�p=
ף�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?              �?      �?        �?wwwwww�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?      �?      �?              �?333333�?�������?              �?      �?              �?        =��<���?�a�a�?      �?        �������?�������?      �?        /�袋.�?F]t�E�?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ1�.hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM/hjh))��}�(h,h/h0M/��h2h3h4hph<�h=Kub������                         x#J@� ��4d�?�           8�@                                  @�~���?|           Ђ@                                   �?>���Rp�?             =@                                  �?ףp=
�?             4@        ������������������������       �                     *@                                    @����X�?             @        ������������������������       �                     @               	                 �(\�?      �?             @        ������������������������       �                     �?        
                        pf�0@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                    @X�<ݚ�?             "@        ������������������������       �                     �?                                   �?      �?              @                                `f�:@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                ���9@�q�q�?             @        ������������������������       �                     �?                                ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               k                    �?�
���?g           �@               h                   �@@x�K��?e             c@              3                     @O����?^             b@               2                    �?�����H�?&             K@              !                     �?(L���?            �E@                                ���;@�q�q�?             @        ������������������������       �                     �?                                 03�=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        "       #                    �?      �?             D@        ������������������������       �                     @        $       -                   �*@؇���X�?            �A@        %       *                 `f�)@����X�?
             ,@       &       )                 `f&'@      �?              @       '       (                   �J@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        +       ,                    :@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        .       1                   �7@���N8�?
             5@        /       0                    ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �        
             &@        4       E                    �?tv?z���?8            �V@        5       @                    �?�E��ӭ�?             B@       6       9                 ���@8�Z$���?             :@        7       8                 �Y�@      �?             @        ������������������������       �                      @        ������������������������       �                      @        :       ?                    �?�C��2(�?             6@        ;       <                   �-@      �?             @        ������������������������       �                     �?        =       >                 �|Y6@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     2@        A       D                    �?���Q��?             $@       B       C                 �|�7@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        F       M                 P�@J��D��?"             K@        G       H                  s@�n_Y�K�?             *@        ������������������������       �                     @        I       L                 �|�9@      �?             $@       J       K                   �2@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        N       ]                 �|�=@��P���?            �D@       O       P                 @33"@ܷ��?��?             =@        ������������������������       �                     $@        Q       X                    �?�S����?             3@        R       S                 Ь�#@�q�q�?             @        ������������������������       �                      @        T       W                 �|�7@      �?             @       U       V                 `F�+@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        Y       \                    �?$�q-�?	             *@       Z       [                   �#@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ^       g                 `f68@      �?             (@       _       b                   &@�q�q�?             "@        `       a                  SE"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        c       f                 03C3@r�q��?             @       d       e                 03�1@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        i       j                      @�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        l       �                    �?�r����?           @z@       m       �                     �?�`�=	�?�            �y@        n       �                    �?�j�'�=�?*            �P@       o       �                   �D@R=6�z�?)            @P@       p       s                 �|�<@�ʻ����?             A@        q       r                 `ffC@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        t                          �@@����"�?             =@       u       z                    �?8����?             7@        v       w                 ���<@�<ݚ�?             "@        ������������������������       �                     @        x       y                 03SA@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        {       |                 `fF<@X�Cc�?             ,@        ������������������������       �                     @        }       ~                   `@@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�q�q�?             @        �       �                   �A@�q�q�?             @        ������������������������       �                     �?        �       �                    C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �B@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �R@��� ��?             ?@       �       �                  �>@ףp=
�?             >@       �       �                 ��>@r�q��?             2@       �       �                   �J@�t����?             1@        �       �                   �G@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @E@�@�9�r�?�            �u@       �       �                    �?����	w�?�            �s@        �       �                    �?�J��%�?            �H@       �       �                 �|Y=@����X�?             E@        �       �                   �5@�\��N��?             3@        �       �                    '@����X�?             @        ������������������������       �                     �?        �       �                 �{@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �9@�q�q�?             (@        ������������������������       �                     @        �       �                  A7@      �?              @       �       �                 �0@r�q��?             @       �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     @���}<S�?             7@        ������������������������       �                     �?        �       �                   @@�C��2(�?             6@       �       �                 ���@r�q��?	             (@       ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �                     $@        �       �                 �y_:@և���X�?             @       �       �                   �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?������?�            �p@        �       �                   `3@@�0�!��?             A@       �       �                 �|Y;@ �Cc}�?             <@        ������������������������       �                     �?        �       �                 ���@�����H�?             ;@        ������������������������       �                     @        �       �                 X��A@R���Q�?             4@       �       �                   @'@�S����?
             3@       ������������������������       �z�G�z�?             .@        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�2@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                   @C@`�q��־?�             m@       �       �                    )@�'B���?�            �k@        �       �                     @z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �@@����Ձ�?�             k@       �       �                    �?@9G��?{            �h@       �       �                     @��R�x��?u            `g@        ������������������������       �                     A@        �       �                   �2@=0�_�?a             c@        �       �                 ��Y @�����H�?             2@        �       �                   �1@      �?              @       �       �                 pf�@r�q��?             @        ������������������������       �                     @        ������������������������       �      �?              @        �       �                 ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �7@`Ӹ����?T            �`@        ������������������������       �                    �D@        �       �                   �;@=QcG��?=            �W@        �       �                 pf� @؇���X�?             5@       �       �                 �Y�@      �?             0@        �       �                 �&b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �:@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 �|�=@���(-�?.            @R@       �       �                 �|Y=@����˵�?&            �M@        ������������������������       �        
             &@        �       �                  sW@      �?             H@        �       �                 pf�@8�Z$���?             *@       ������������������������       �                      @        ������������������������       ����Q��?             @        �       �                 ��) @��?^�k�?            �A@       ������������������������       �                     ;@        �       �                 pf� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     "@        �       �                   @A@�����?             5@        �       �                     @����X�?             @        �       �                    1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        �       �                     @���|���?             &@        �       �                    4@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 pf� @      �?              @       �       �                   �C@���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     >@        ������������������������       �                      @              &                    �? ��?�?F            @[@                                �?�+I�9��?<            @V@                             ���P@HP�s��?3            �R@                              `�>P@�㙢�c�?             7@                                5@�����?             5@                              `f�K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        	      
                p��K@�}�+r��?             3@        ������������������������       �                     &@                              �5L@      �?              @                                @F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                 �? ��WV�?#             J@       ������������������������       �                    �E@                                 �?�<ݚ�?             "@                                �?����X�?             @                              �	U@���Q��?             @        ������������������������       �                     �?                              �|Y;@      �?             @        ������������������������       �                      @                              0�c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @              %                  �G@����X�?	             ,@                              �(\�?�θ�?             *@        ������������������������       �                     @        !      "                   $@�q�q�?             "@        ������������������������       �                      @        #      $                   �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        '      *                   �?z�G�z�?
             4@        (      )                    @�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        +      ,                    @���!pc�?             &@        ������������������������       �                      @        -      .                   ;@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M/KK��h2h3h4hVh<�h=Kub��������������`uv��?,J>��?�� [	��?�L�I�-�?GX�i���?�i��F�?�������?�������?              �?�$I�$I�?�m۶m��?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        r�q��?�q�q�?              �?      �?      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?!�G˭�?�#pi��?�?ssssss�?�8��8��?��8��8�?�q�q�?�q�q�?w�qG��?⎸#��?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?              �?�$I�$I�?۶m۶m�?�$I�$I�?�m۶m��?      �?      �?�$I�$I�?�m۶m��?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�a�a�?��y��y�?      �?      �?      �?                      �?              �?              �?a�`��??�>��?r�q��?�q�q�?;�;��?;�;��?      �?      �?              �?      �?        F]t�E�?]t�E�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?�������?      �?      �?      �?                      �?      �?        �^B{	��?_B{	�%�?ى�؉��?;�;��?              �?      �?      �?�$I�$I�?�m۶m��?      �?                      �?      �?        ������?�����?��=���?a���{�?      �?        (������?^Cy�5�?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�؉�؉�?;�;��?�q�q�?�q�q�?              �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        9��8���?�q�q�?              �?      �?        �������?�?��6���?�H%�e�?�&�l���?m��&�l�?Wj�Vj��?S+�R+��?�������?<<<<<<�?�������?�������?              �?      �?        	�=����?�i��F�?d!Y�B�?8��Moz�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        %I�$I��?�m۶m��?      �?        �q�q�?r�q��?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �{����?�B!��?�������?�������?�������?UUUUUU�?<<<<<<�?�?      �?      �?      �?                      �?      �?                      �?      �?                      �?      �?        �}����?�DZ/`�?��td�@�?�Z܄��?c}h���?9/����?�m۶m��?�$I�$I�?�5��P�?y�5���?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?                      �?�������?�������?      �?              �?      �?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?        ӛ���7�?d!Y�B�?      �?        ]t�E�?F]t�E�?�������?UUUUUU�?      �?        333333�?�������?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?        ؽ�u�{�?B�P�"�?ZZZZZZ�?�������?%I�$I��?۶m۶m�?      �?        �q�q�?�q�q�?      �?        333333�?333333�?(������?^Cy�5�?�������?�������?      �?              �?              �?      �?      �?                      �?��6���?r؃H{�?��$j�?镱��^�?�������?�������?      �?                      �?��}��?�`^0/��?������?9/���?��rD���?�и[�?      �?        ��S��S�?p�pŪ?�q�q�?�q�q�?      �?      �?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?                      �?      �?        ?�>��?l�l��?      �?        x6�;��?AL� &W�?۶m۶m�?�$I�$I�?      �?      �?�������?�������?      �?                      �?      �?        333333�?�������?      �?                      �?��իW��?�P�B�
�?W'u_�?��/���?      �?              �?      �?;�;��?;�;��?      �?        333333�?�������?_�_��?�A�A�?      �?              �?      �?              �?      �?              �?              �?        =��<���?�a�a�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?333333�?�������?UUUUUU�?UUUUUU�?      �?              �?              �?              �?        ���]8��?߅���]�?�as�ü?�3��g�?{�G�z�?q=
ףp�?d!Y�B�?�7��Mo�?�a�a�?=��<���?      �?      �?      �?                      �?(�����?�5��P�?              �?      �?      �?      �?      �?              �?      �?                      �?      �?        ;�;��?O��N���?              �?�q�q�?9��8���?�$I�$I�?�m۶m��?�������?333333�?      �?              �?      �?              �?      �?      �?              �?      �?                      �?              �?�$I�$I�?�m۶m��?�؉�؉�?ى�؉��?              �?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?        �������?�������?�q�q�?�q�q�?              �?      �?        F]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg�)hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM!hjh))��}�(h,h/h0M!��h2h3h4hph<�h=Kub������       h                    �?���?Y��?�           8�@               #                    �?�����?�             q@               "                    @8��8���?>             X@                                  �?��E�B��?=            �W@                               `�@1@������?.            �Q@                                    @X�<ݚ�?             2@        ������������������������       �                     @                                   �?և���X�?
             ,@       	       
                   �,@      �?             $@        ������������������������       �                      @                                �%@      �?              @        ������������������������       �                     �?                                  �-@����X�?             @        ������������������������       �                     @                                ���,@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   �?      �?             @        ������������������������       �                      @                                �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �H@ pƵHP�?!             J@       ������������������������       �                     D@                                ���I@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@                                    @      �?             8@        ������������������������       �                     @               !                    �?R���Q�?             4@                                �&�@�KM�]�?             3@        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     �?        ������������������������       �                      @        $       /                    !@�z/sT�?j            @f@        %       &                    �?�����?             5@        ������������������������       �                     @        '       *                 �̌5@�r����?
             .@        (       )                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        +       ,                 03�=@$�q-�?             *@       ������������������������       �                     @        -       .                 ��T?@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        0       c                    @�(T���?_            �c@       1       2                    (@�SW���?Y            �b@        ������������������������       �                     $@        3       D                     @�-١�:�?T            @a@       4       C                    �?Pq�����?5            @U@       5       :                   �B@Hm_!'1�?             �H@       6       9                   �7@��?^�k�?            �A@        7       8                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ;@        ;       <                     �?d}h���?
             ,@        ������������������������       �                     @        =       >                   �C@�z�G��?             $@        ������������������������       �                      @        ?       @                    5@      �?              @       ������������������������       �                     @        A       B                   �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     B@        E       N                   �7@l`N���?            �J@        F       K                    �?j���� �?             1@       G       H                   �2@�eP*L��?             &@        ������������������������       �                     @        I       J                 8�!@      �?              @       ������������������������       �                     @        ������������������������       �                      @        L       M                 ���5@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        O       T                   �:@�q�q�?             B@        P       Q                   �9@$�q-�?             *@       ������������������������       �                      @        R       S                 xF�'@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        U       b                   @B@
;&����?             7@       V       _                    �?�G��l��?             5@       W       X                 �|�<@���Q��?             .@        ������������������������       �                     �?        Y       Z                 pf�$@X�Cc�?             ,@        ������������������������       �                     @        [       \                   �>@ףp=
�?             $@       ������������������������       �                     @        ]       ^                 03�1@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        `       a                 ���5@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        d       e                    @�����H�?             "@        ������������������������       �                     @        f       g                   @C@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        i       v                    @b������?           P{@        j       s                    �?     ��?             0@       k       l                 �G�?"pc�
�?             &@        ������������������������       �                     @        m       n                 03�6@���Q��?             @        ������������������������       �                      @        o       p                   A@�q�q�?             @        ������������������������       �                     �?        q       r                     @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        t       u                     @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        w       �                 ��K.@�]C9��?           Pz@       x       �                     @Dg�-N�?�            q@        y       |                    4@$�q-�?)            @P@        z       {                    &@�<ݚ�?             "@        ������������������������       ��q�q�?             @        ������������������������       �                     @        }       ~                     �?�h����?$             L@        ������������������������       �                     @               �                   �)@0G���ջ?"             J@        ������������������������       �                     8@        �       �                    �? �Cc}�?             <@        ������������������������       �                     @        �       �                 �|Y<@H%u��?             9@        ������������������������       �                     "@        �       �                 �|�=@     ��?             0@        ������������������������       �                     �?        �       �                   �*@�r����?             .@       �       �                    @@�<ݚ�?             "@        ������������������������       �                      @        �       �                   �A@����X�?             @        ������������������������       �                     �?        �       �                   @D@r�q��?             @        ������������������������       �                      @        �       �                    G@      �?             @       ������������������������       �      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���@ȵHPS!�?�             j@        ������������������������       �                     9@        �       �                   �0@(��+�?y            �f@        �       �                 �Yu$@      �?             @       �       �                 pFD!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @@@x疑��?v            `f@       �       �                   �>@�npº��?f            �b@       �       �                 ��@L�
�$�?a            �a@        ������������������������       �                      @        �       �                    �?��27
��?`            `a@        �       �                    �?tk~X��?             B@       �       �                    8@�q�q�?             8@        ������������������������       �                     @        �       �                 ���@�����?             5@        ������������������������       �                     @        �       �                   �<@؇���X�?             ,@        ������������������������       �                     @        �       �                 �|Y=@z�G�z�?             $@        ������������������������       �                     �?        �       �                 �|�=@�����H�?             "@       �       �                   @@      �?              @       ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                  ��@r�q��?
             (@        ������������������������       �                     @        ������������������������       �      �?              @        �       �                   �2@�b�E�V�?E            �Y@        �       �                   �1@�q�q�?             @        ������������������������       �                     @        �       �                 ��Y @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �:@�*v��?A            @X@        �       �                 @3�@��Y��]�?            �D@       ������������������������       �                     =@        �       �                    4@�8��8��?             (@        �       �                 `�8"@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ��) @4և����?"             L@       �       �                 �&B@�?�|�?            �B@        �       �                 pf�@�����H�?             "@       ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     <@        �       �                   �;@���y4F�?	             3@        ������������������������       �                     �?        �       �                 pf� @r�q��?             2@        ������������������������       �                     @        ������������������������       �                     .@        �       �                   �@���Q��?             $@        ������������������������       �                     �?        �       �                 �?�@�q�q�?             "@        ������������������������       �                     @        �       �                   �?@      �?             @        ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     <@        �                         @C@���+�?]            �b@       �       �                 �y�/@�ԇ���?C            �Y@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 `fFJ@.��Zr��??            @X@       �       �                     �?����>�?0            �R@        �       �                    �?�99lMt�?            �C@       �       �                   �;@؀�:M�?            �B@        ������������������������       �                     @        �       �                   �>@�!���?             A@        �       �                 X�,@@j���� �?	             1@       �       �                    �?      �?             ,@        �       �                 �ܵ<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @>@      �?             (@       �       �                 ��<:@      �?              @        ������������������������       �                     @        �       �                 `fF<@���Q��?             @       �       �                 �|�<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �|�<@�IєX�?             1@        �       �                 `f�D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             *@        ������������������������       �                      @        �       �                    #@b�h�d.�?            �A@        �       �                 03�8@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�r����?             >@        �       �                     @X�<ݚ�?             "@        ������������������������       �                     @        �       �                 03�7@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        �                          �?
;&����?             7@       �                          �?�G��l��?             5@        �       �                 p"4W@�q�q�?             @        ������������������������       �                     �?                                  �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?                                �7@���Q��?
             .@        ������������������������       �                      @                                   @�	j*D�?             *@                                �?�q�q�?             "@             
                `f�K@؇���X�?             @              	                   @@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                 >@      �?             @                                ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                               x;K@�r����?            �F@                                 �?�FVQ&�?            �@@                                �H@      �?	             0@        ������������������������       �                      @                                 K@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             1@                              0��M@�q�q�?             (@        ������������������������       �                      @                                 @H@z�G�z�?             $@                                �G@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M!KK��h2h3h4hVh<�h=Kub��������������� 3��?@Bx���?������?����?�������?UUUUUU�?AL� &W�?�l�w6��?PuPu�?,��+���?�q�q�?r�q��?              �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?              �?      �?              �?      �?        ;�;��?'vb'vb�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?333333�?333333�?(�����?�k(���?      �?                      �?      �?              �?        <��x��?bs���?�a�a�?=��<���?              �?�?�������?      �?      �?              �?      �?        ;�;��?�؉�؉�?              �?�$I�$I�?۶m۶m�?      �?                      �?F����?�\�:�2�?Z7�"�u�?S�n0E�?      �?        s��\;�?~F��Q��?�?~~~~~~�?9/���?Y�Cc�?�A�A�?_�_��?      �?      �?      �?                      �?              �?۶m۶m�?I�$I�$�?              �?333333�?ffffff�?      �?              �?      �?              �?      �?      �?              �?      �?                      �?�R���?
�[���?ZZZZZZ�?�������?]t�E�?t�E]t�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?�؉�؉�?;�;��?      �?        �������?�������?              �?      �?        Y�B��?�Mozӛ�?��y��y�?1�0��?�������?333333�?      �?        �m۶m��?%I�$I��?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �q�q�?�q�q�?      �?        �������?�������?              �?      �?        �eJV��?Fh֊���?      �?      �?F]t�E�?/�袋.�?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?�������?              �?      �?        �-шs��?�I��1��?�ə�ə�?�1�1�?�؉�؉�?;�;��?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?        vb'vb'�?�؉�؉�?      �?        %I�$I��?۶m۶m�?      �?        )\���(�?���Q��?      �?              �?      �?              �?�������?�?9��8���?�q�q�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?              �?        ��N��N�?�؉�؉�?      �?        q�����?;ڼOq��?      �?      �?      �?      �?              �?      �?                      �?��fh�>�?59ȼ��?�2n���?�4G�#��?qJ��O$�?{�e�ݾ?              �?�j����?p�l�:��?r�q��?9��8���?UUUUUU�?�������?              �?=��<���?�a�a�?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?�q�q�?�q�q�?      �?      �?      �?      �?      �?              �?        �������?UUUUUU�?      �?              �?      �?�jch���?��,�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���AG�? tT����?8��18�?������?      �?        UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?      �?      �?              �?        I�$I�$�?�m۶m۶?*�Y7�"�?к����?�q�q�?�q�q�?      �?              �?      �?      �?        6��P^C�?(������?              �?�������?UUUUUU�?              �?      �?        333333�?�������?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?      �?      �?        �n0E>��?�"�u�)�?�`�����?#>�Tr^�?UUUUUU�?�������?              �?      �?        �:*���?T���t�?�u�)�Y�?���L�?5H�4H��?�o��o��?E>�S��?v�)�Y7�?              �?�������?�������?ZZZZZZ�?�������?      �?      �?      �?      �?      �?                      �?      �?      �?      �?      �?      �?        333333�?�������?      �?      �?              �?      �?              �?                      �?              �?�?�?      �?      �?              �?      �?              �?              �?        ;��:���?_�_��?333333�?�������?              �?      �?        �������?�?r�q��?�q�q�?      �?        �������?�������?              �?      �?              �?        Y�B��?�Mozӛ�?��y��y�?1�0��?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?�������?333333�?      �?        ;�;��?vb'vb'�?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?      �?      �?              �?      �?                      �?      �?        �������?�?>����?|���?      �?      �?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�]_AhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       n                    �?^����[�?�           8�@               _                 ��T?@H��0~��?�            �o@              ^                    @ҐϿ<��?k            �f@                                  (@��Ж�H�?j            `f@                                   �?l��[B��?             =@                                `��+@d}h���?             ,@        ������������������������       �                     @                                   �?      �?              @        	       
                 `�@1@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                   @      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                   !@z�G�z�?             .@                                   @      �?              @                               `f�:@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @               3                     @�M;q��?Z            �b@               .                 03;<@\#r��?%            �N@                                 �&@�NW���?!            �J@                                  �J@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?               #                   @4@=QcG��?            �G@               "                   �*@ 7���B�?             ;@                                  �?�IєX�?             1@        ������������������������       �                     �?                !                    B@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �                     $@        $       %                     �?ףp=
�?             4@        ������������������������       �                     @        &       )                   �;@      �?             0@        '       (                   �9@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        *       +                   �E@�8��8��?	             (@       ������������������������       �                      @        ,       -                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        /       2                     �?      �?              @        0       1                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        4       5                   �1@�L��7Q�?5            @V@        ������������������������       �                      @        6       C                    �?L����?0            @T@        7       >                 �YU&@R�}e�.�?             :@       8       =                    �?r�q��?             2@       9       <                 ���@�t����?
             1@        :       ;                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     �?        ?       @                    5@      �?              @        ������������������������       �                     �?        A       B                 ��.@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        D       E                  s@ؓ��M{�?            �K@        ������������������������       �                     @        F       W                   �>@x�K��?            �I@       G       V                   �;@�����?             C@       H       I                 ���@��
ц��?             :@        ������������������������       �                     @        J       K                 �&B@�û��|�?             7@        ������������������������       �                     @        L       U                    �?�G�z��?             4@       M       R                   �9@������?
             .@       N       Q                   �4@�����H�?             "@        O       P                   �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        S       T                 pf(@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        X       ]                    �?�n_Y�K�?             *@       Y       \                   @D@�eP*L��?             &@       Z       [                 03�1@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        `       i                 ��R@�X�<ݺ?-             R@        a       b                    �? �Cc}�?             <@        ������������������������       �                     $@        c       f                 �|Y?@r�q��?             2@        d       e                 @3cN@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        g       h                    @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        j       k                    �?`���i��?             F@       ������������������������       �                    �C@        l       m                    '@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        o       ~                    '@�i����?!           �|@        p       q                     @�+e�X�?             9@        ������������������������       �                      @        r       s                    �?ҳ�wY;�?             1@        ������������������������       �                     �?        t       u                    @     ��?
             0@        ������������������������       �                     @        v       }                 pf�C@8�Z$���?             *@       w       x                    �?�8��8��?             (@        ������������������������       �                     @        y       z                 `f�9@؇���X�?             @        ������������������������       �                     @        {       |                 ��T?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?               �                    �?�؏�9�?           �z@        �       �                   �;@x�(�3��?1            @S@        �       �                      @�q�q�?             8@        �       �                  �}S@�	j*D�?             *@        ������������������������       �                     @        �       �                   �1@և���X�?             @        ������������������������       �                      @        �       �                   �8@z�G�z�?             @        ������������������������       �                     @        �       �                    :@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��y@�eP*L��?             &@        ������������������������       �                      @        �       �                 H�%@X�<ݚ�?             "@       �       �                    �?�q�q�?             @       �       �                   �7@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     �?�iʫ{�?"            �J@        �       �                  xCH@      �?             8@       �       �                 �|�=@�8��8��?             (@        �       �                 ��2>@r�q��?             @        �       �                 �ܵ<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�q�q�?             (@       �       �                 @��V@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                 �w�q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��,@ܷ��?��?             =@       ������������������������       �                     7@        �       �                 �|�=@      �?             @       �       �                     @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ��D:@��g�g�?�             v@       �       �                   �2@�E�J��?�            �p@        �       �                 ��Y @������?             1@        �       �                   �1@���Q��?             $@       �       �                 pf�@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @        �       �                  s@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?$Q�q�?�            �o@        �       �                 X��A@�IєX�?             A@       �       �                   `3@ 	��p�?             =@       ������������������������       �                     :@        �       �                 03�7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|�=@HQ˄�ľ?�            @k@       �       �                    �?�d����?a            @a@       �       �                   �;@�?�0�!�?_             a@       �       �                     @      �?8             T@        �       �                    4@@4և���?             ,@        ������������������������       �      �?              @        ������������������������       �        
             (@        �       �                   �:@�FVQ&�?,            �P@       �       �                 ���@     �?*             P@        �       �                 ���@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        �       �                   @4@�O4R���?#            �J@        �       �                   �3@�8��8��?             (@       ������������������������       �                     @        �       �                 @3�@z�G�z�?             @        �       �                 P�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@        �       �                 �� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        '             L@        ������������������������       �                      @        �       �                   �*@���(\��?/             T@       �       �                   @A@R���Q�?"             N@        �       �                   �@@�z�G��?             >@       �       �                   @@@�+e�X�?             9@       �       �                    $@����X�?             5@       �       �                 �̌!@      �?             (@       �       �                   �>@���Q��?             $@        ������������������������       �                      @        �       �                   �?@      �?              @        ������������������������       �                     �?        �       �                 P�@և���X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       ����Q��?             @        ������������������������       �                     >@        ������������������������       �                     4@        �                           �?�t����?2            @U@       �                          �?ҳ�wY;�?(             Q@       �                          �>@���@M^�?$             O@        �       �                   �J@
j*D>�?             :@       �       �                 `f�;@�����?	             3@       �       �                 X�,@@ףp=
�?             $@        �       �                 �|�<@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 X��B@X�<ݚ�?             "@       �       �                 �|Y=@�q�q�?             @       �       �                   @>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    R@����X�?             @       ������������������������       �                     @        ������������������������       �                      @                                @H@      �?             B@                               �E@z�G�z�?             >@                             �|Y>@�q�q�?             2@                             �|�<@r�q��?             (@                              `f�D@�q�q�?             @        ������������������������       �                     �?                              ��I@z�G�z�?             @        ������������������������       �                      @        	      
                   7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                               x#J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@                              ���T@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                              0�H@�IєX�?
             1@        ������������������������       �                     $@                              �|�>@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������C�B���?�x�z���?�������?�������?mާ�d�?������?k��P�?J���s�?���=��?GX�i���?۶m۶m�?I�$I�$�?              �?      �?      �?      �?      �?      �?                      �?      �?      �?              �?      �?        �������?�������?      �?      �?�������?UUUUUU�?              �?      �?                      �?      �?        ƒ_,���?�6�i��?XG��).�?��:��?�x+�R�?萚`���?UUUUUU�?�������?              �?      �?        AL� &W�?x6�;��?h/�����?	�%����?�?�?              �?      �?      �?              �?      �?                      �?�������?�������?              �?      �?      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?��MmjS�?%+Y�JV�?              �?�5?,R�?#e�����?�;�;�?'vb'vb�?UUUUUU�?�������?�?<<<<<<�?�������?333333�?              �?      �?                      �?      �?              �?      �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?	� O	�?�־a��?              �?ssssss�?�?Q^Cy��?^Cy�5�?�;�;�?�؉�؉�?              �?8��Moz�?��,d!�?      �?        �������?�������?wwwwww�?�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?                      �?      �?        ى�؉��?;�;��?]t�E�?t�E]t�?      �?      �?              �?      �?              �?                      �?      �?        �q�q�?��8��8�?۶m۶m�?%I�$I��?              �?UUUUUU�?�������?�$I�$I�?�m۶m��?              �?      �?        F]t�E�?]t�E�?              �?      �?        F]t�E�?F]t�E�?              �?�������?�������?      �?                      �?Q^Cy��?����k�?���Q��?R���Q�?              �?�������?�������?      �?              �?      �?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ^�Ԇ��?�Bp��1�?(�Y�	q�?�wL��?�������?�������?;�;��?vb'vb'�?              �?�$I�$I�?۶m۶m�?              �?�������?�������?      �?              �?      �?              �?      �?        t�E]t�?]t�E�?      �?        �q�q�?r�q��?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        
�[���?�琚`��?      �?      �?UUUUUU�?UUUUUU�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?333333�?�������?              �?      �?              �?      �?      �?                      �?��=���?a���{�?      �?              �?      �?      �?      �?      �?                      �?      �?        ي����?��}ylE�?�-���?��~���?xxxxxx�?�?333333�?�������?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        ~��}���?AA�?�?�?������?�{a���?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ߅����?��p�?��\;0��?)�3J���?�������?�����Ң?      �?      �?n۶m۶�?�$I�$I�?      �?      �?      �?        >����?|���?     ��?      �?/�袋.�?F]t�E�?      �?                      �?:�&oe�?�x+�R�?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?      �?      �?                      �?      �?              �?              �?      �?      �?                      �?      �?              �?        ffffff�?�����̼?333333�?333333�?ffffff�?333333�?R���Q�?���Q��?�m۶m��?�$I�$I�?      �?      �?333333�?�������?      �?              �?      �?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?333333�?      �?              �?        �������?�������?�������?�������?�s�9��?�c�1��?;�;��?b'vb'v�?^Cy�5�?Q^Cy��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?r�q��?�q�q�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �m۶m��?�$I�$I�?      �?                      �?      �?      �?�������?�������?UUUUUU�?UUUUUU�?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?      �?        �?�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJL�OhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       @                    �?�E	�rQ�?�           8�@                                    @�YP-��?�            `o@                                 @L@pJQg���?S            �`@                                  �? �|ك�?O            �^@                                  �H@�(\����?             D@       ������������������������       �                    �B@               
                   �J@�q�q�?             @              	                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        6            �T@                                `f�2@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @               1                 @�+@�m����?O            �]@                                 �3@r֛w���?+             O@        ������������������������       �                     5@               0                    A@hP�vCu�?            �D@              %                 �̌@�99lMt�?            �C@              $                    �?��2(&�?             6@                               pff@�����?             5@                                   �?�q�q�?             @        ������������������������       �                     �?                                �|�9@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?�X�<ݺ?             2@       ������������������������       �                     &@                                ���@؇���X�?             @        ������������������������       �                     �?                #                 �&B@r�q��?             @       !       "                   �7@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        &       /                 ��&@ҳ�wY;�?             1@       '       .                 `��!@d}h���?
             ,@        (       )                 �?�@      �?             @        ������������������������       �                     �?        *       -                 ��� @���Q��?             @       +       ,                   �9@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        2       ;                 ��*4@      �?$             L@        3       4                    @     ��?             @@        ������������������������       �                     @        5       6                 ��.@��X��?             <@        ������������������������       �                     .@        7       8                 ���1@�	j*D�?	             *@       ������������������������       �                      @        9       :                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        <       =                 ��T?@ �q�q�?             8@       ������������������������       �                     0@        >       ?                    @      �?              @       ������������������������       �                     @        ������������������������       �                     �?        A       x                    �?Xf1�
�?,           �|@        B       a                     �?�	j*D�?5            �S@        C       `                    �?���Q��?            �A@       D       Y                   @F@4���C�?            �@@       E       R                 �D�G@��Q��?             4@       F       Q                    C@�eP*L��?             &@       G       H                 �|�;@�q�q�?             "@        ������������������������       �                     �?        I       P                   �A@      �?              @       J       O                   @@@�q�q�?             @       K       N                 �|�=@z�G�z�?             @       L       M                 ��2>@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        S       T                 ��)e@�����H�?             "@       ������������������������       �                     @        U       V                    �?      �?             @        ������������������������       �                     �?        W       X                    >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Z       _                    �?$�q-�?	             *@       [       \                 xSQ@�����H�?             "@       ������������������������       �                     @        ]       ^                   �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        b       q                    �?>��C��?            �E@       c       p                 �|Y=@@�0�!��?             A@        d       e                    5@և���X�?	             ,@        ������������������������       �                     @        f       o                  A7@���Q��?             $@       g       h                   �6@�q�q�?             "@        ������������������������       �                     @        i       j                   @@      �?             @        ������������������������       �                      @        k       n                 �0@      �?             @       l       m                    <@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@        r       s                 ��y&@X�<ݚ�?             "@        ������������������������       �                     @        t       w                 �|Y;@�q�q�?             @        u       v                 pV�C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        y       �                    @���Jh��?�            �w@        z                          �;@������?             .@       {       ~                    @ףp=
�?             $@        |       }                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��T?@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                     �?0<o�Ɲ�?�            �v@        �       �                    �?8^s]e�?$             M@       �       �                    R@��X��?"             L@       �       �                  i?@l��
I��?!             K@       �       �                    K@      �?             8@       �       �                 03:@�q�q�?             2@        ������������������������       �                     @        �       �                   �F@z�G�z�?             .@       �       �                 �|�?@ףp=
�?             $@       �       �                 �|�<@z�G�z�?             @        ������������������������       �                      @        �       �                 `fF<@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   `G@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 03�U@�r����?             >@       �       �                    A@@4և���?             <@        �       �                   �;@����X�?             @        �       �                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y>@z�G�z�?             @       ������������������������       �                     @        �       �                 0��J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                     @�luL3�?�            Ps@        �       �                    4@$�q-�?%             J@        �       �                   �1@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 �|�=@ �q�q�?#             H@        �       �                    �?�C��2(�?             6@       �       �                 �|Y=@�����?             5@       ������������������������       �        
             1@        �       �                    @      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     :@        �       �                 �T�I@�pe��?�            p@       �       �                  ��@����y7�?�            @o@        �       �                   �8@@��8��?             H@        �       �                    7@��S�ۿ?             .@       ������������������������       �                     $@        �       �                 `fF@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �@@        �       �                    �?x�7Fb��?�            @i@       �       �                    �?�+�$f��?~            �h@        �       �                   �2@�n`���?             ?@        ������������������������       �                     @        �       �                    �?�<ݚ�?             ;@       �       �                 �|Y=@�θ�?             :@        ������������������������       �                      @        �       �                 X��A@r�q��?             8@       �       �                 ��(@"pc�
�?             6@       ������������������������       �������?             1@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?|T(W�j�?l            �d@       �       �                   �4@�d	���?f            �c@        �       �                 ��Y @�<ݚ�?             B@       �       �                 �?�@���Q��?             4@        ������������������������       �                      @        �       �                 @3�@�q�q�?             (@        ������������������������       ��q�q�?             @        �       �                   �3@�q�q�?             "@       �       �                   �2@      �?              @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     0@        �       �                   �>@ @|���?N            �^@       �       �                 �?$@P��BNֱ?3            �T@        �       �                 �|�;@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        �       �                 ��) @pY���D�?0            �S@       ������������������������       �        !             M@        �       �                   �:@�����?             5@        ������������������������       �                     @        �       �                   �;@�r����?
             .@        ������������������������       �                     �?        �       �                 �|Y=@@4և���?	             ,@        ������������������������       �                     @        �       �                 pf� @ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �?@��-�=��?            �C@        ������������������������       �                      @        �       �                   @@@@-�_ .�?            �B@        �       �                 ��I @؇���X�?             @       �       �                 �?�@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        �       �                 @3�@(;L]n�?             >@        �       �                   @C@ףp=
�?             $@        ������������������������       �                     @        �       �                 �?�@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �       �                    0@؇���X�?             @        �       �                   �5@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    $@r�q��?             @        �       �                 83�@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                       p�O@և���X�?             @                              �|�>@      �?             @                                ;@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������JP���?7j_Q��?(;r���?6q�9�?�qA��?s���7G�?�h
���?�_��e��?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?�������?�������?      �?                      �?�V'u�?��}ylE�?�B!��?���{��?              �?������?��18��?�o��o��?5H�4H��?t�E]t�?��.���?�a�a�?=��<���?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �q�q�?��8��8�?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?�������?�������?              �?      �?                      �?      �?        �������?�������?I�$I�$�?۶m۶m�?      �?      �?      �?        �������?333333�?      �?      �?      �?                      �?              �?      �?                      �?      �?              �?      �?      �?      �?              �?n۶m۶�?%I�$I��?      �?        ;�;��?vb'vb'�?              �?�������?�������?              �?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?���(�?vI�ø_�?vb'vb'�?;�;��?333333�?�������?m��&�l�?'�l��&�?ffffff�?�������?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?              �?                      �?      �?                      �?�q�q�?�q�q�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�؉�؉�?;�;��?�q�q�?�q�q�?      �?              �?      �?              �?      �?              �?              �?        $�;��?qG�w��?ZZZZZZ�?�������?�$I�$I�?۶m۶m�?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?      �?      �?                      �?              �?      �?              �?        r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?�&�eL��?�d�h��?�?wwwwww�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?�������?      �?                      �?���>��?%e��?|a���?	�=����?n۶m۶�?%I�$I��?Lh/����?h/�����?      �?      �?UUUUUU�?UUUUUU�?      �?        �������?�������?�������?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?333333�?      �?                      �?      �?        �������?�?n۶m۶�?�$I�$I�?�m۶m��?�$I�$I�?      �?      �?      �?                      �?�������?�������?      �?              �?      �?      �?                      �?      �?                      �?              �?      �?        �+&��?NZ�Ϯ�?�؉�؉�?;�;��?      �?      �?      �?                      �?�������?UUUUUU�?]t�E�?F]t�E�?=��<���?�a�a�?      �?              �?      �?      �?                      �?      �?              �?        ]�\�\��?���?!�rh���?�~j�t��?UUUUUU�?UUUUUU�?�������?�?      �?        �������?�������?              �?      �?              �?        �<�]?[�?Y�&�?�Cc}h�?/�����?�9�s��?�c�1��?      �?        9��8���?�q�q�?ى�؉��?�؉�؉�?              �?�������?UUUUUU�?/�袋.�?F]t�E�?xxxxxx�?�?      �?              �?              �?        ��YΟ��?�0�Ӹ?��JG��?�0���M�?9��8���?�q�q�?333333�?�������?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?        "XG��)�?�}�K�`�?��FS���?���ˊ��?      �?      �?      �?        UUUUUU�?UUUUUU�?a~W��0�?�3���?      �?        =��<���?�a�a�?      �?        �������?�?              �?n۶m۶�?�$I�$I�?      �?        �������?�������?              �?      �?        }˷|˷�?�A�A�?              �?S�n0E�?к����?۶m۶m�?�$I�$I�?�������?�������?      �?              �?      �?      �?        �������?�?�������?�������?      �?        �������?�������?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        �������?UUUUUU�?      �?      �?              �?      �?              �?        �$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��lhG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiM%hjh))��}�(h,h/h0M%��h2h3h4hph<�h=Kub������       �                 `�X.@>AU`�z�?�           8�@                                  /@�+e�X�?�            pw@               
                    �?�t����?             1@               	                    �?�<ݚ�?             "@                                 �,@�q�q�?             @        ������������������������       �                     @                                  �-@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @               ?                    �?4F娥2�?�            `v@                                   �9@�sly47�?3            �R@                                  �6@X�<ݚ�?             ;@                               �[$@�d�����?             3@                                  �?@�0�!��?             1@        ������������������������       �                     @                                   4@�θ�?             *@                                  �?"pc�
�?             &@                               �&B@�<ݚ�?             "@                                P��@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                ��y!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                pf�@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        !       >                 �B,@�q�q��?              H@       "       +                    �?:	��ʵ�?            �F@        #       $                     @ףp=
�?             4@        ������������������������       �                     @        %       (                 ���@�t����?             1@        &       '                 �Y�@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        )       *                    �?@4և���?	             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ,       -                   �;@�+e�X�?             9@        ������������������������       �                     "@        .       5                 `f�$@      �?             0@        /       4                    �?r�q��?             @       0       1                 �|Y>@z�G�z�?             @        ������������������������       �                     @        2       3                  SE"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        6       7                   �'@ףp=
�?             $@        ������������������������       �                     �?        8       9                   �B@�����H�?             "@       ������������������������       �                     @        :       =                   �*@      �?             @       ;       <                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        @       U                     @��|C_�?�            �q@        A       B                     �?�����H�?"             K@        ������������������������       �                     @        C       T                   @A@�t����?             �I@       D       K                 `fF)@r�q��?             B@        E       J                    &@�����H�?
             2@       F       G                    @8�Z$���?             *@        ������������������������       �                     �?        H       I                    5@r�q��?             (@        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     @        L       S                    @@�<ݚ�?             2@       M       N                 �|Y;@�r����?	             .@       ������������������������       �                     @        O       R                 �|�=@      �?              @       P       Q                 ��,@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       ��q�q�?             @        ������������������������       �                     .@        V       �                    �?T�����?�            �l@       W       �                 ���"@$�q-�?�            �k@       X       g                    �? "��u�?~             i@        Y       Z                 ���@�>����?!             K@        ������������������������       �        
             0@        [       ^                 ���@�KM�]�?             C@        \       ]                 �|�=@���Q��?             @       ������������������������       �      �?             @        ������������������������       �                     �?        _       f                 P�J@�FVQ&�?            �@@       `       a                  ��@�C��2(�?             6@        ������������������������       �                     @        b       c                 �|Y=@�t����?             1@        ������������������������       �                     �?        d       e                 X��A@      �?
             0@       ������������������������       ��8��8��?             (@        ������������������������       �                     @        ������������������������       �                     &@        h       o                   �3@F��}��?]            @b@        i       j                   �2@�����H�?             2@       ������������������������       �        
             &@        k       l                 �?�@����X�?             @       ������������������������       �                     @        m       n                 0S5 @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        p       q                 ���@     �?N             `@        ������������������������       �        	             4@        r       s                   �7@�X�<ݺ?E             [@        ������������������������       �                     <@        t       u                 ���@��(\���?7             T@        ������������������������       �                      @        v       }                 �?�@�7��?6            �S@       w       |                 �?$@`���i��?             F@        x       {                 �|Y>@��S�ۿ?             .@       y       z                 ���@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     =@        ~       �                 @3�@l��\��?             A@               �                   �A@�q�q�?             @       �       �                    >@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?        �       �                 ��) @h�����?             <@       ������������������������       �                     3@        �       �                 �|�>@�����H�?             "@        �       �                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    <@���N8�?             5@        ������������������������       �                     "@        �       �                    (@�q�q�?             (@        �       �                   �?@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                  x#J@��Bu��?�             u@       �       �                    �?�6)��?�            �k@       �       �                    �?���Q��?U            @`@        �       �                 ��4=@��Q��?             4@        ������������������������       �                     @        �       �                     �?j���� �?             1@       �       �                    �?     ��?             0@        ������������������������       �                     @        �       �                    H@�	j*D�?
             *@       �       �                  Y>@      �?              @        ������������������������       �                     @        �       �                    C@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?8�A�0��?E            �[@        �       �                   �;@"pc�
�?            �@@        �       �                   �7@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�>����?             ;@        ������������������������       �                     @        �       �                   �E@���}<S�?             7@       ������������������������       �        	             0@        �       �                   @G@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �J@N��c��?1            @S@       �       �                   �H@���!pc�?*            �P@       �       �                     �?���N8�?(            �O@        �       �                    D@4���C�?            �@@       �       �                   @@@��
ц��?             :@       �       �                   �;@���Q��?             4@        ������������������������       �                     @        �       �                   �>@      �?             0@        �       �                 ��<:@և���X�?             @        ������������������������       �                     �?        �       �                   @>@�q�q�?             @       �       �                 `fF<@���Q��?             @        �       �                 �|�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @        �       �                     @(;L]n�?             >@        ������������������������       �        	             .@        �       �                 �|�:@��S�ۿ?             .@        ������������������������       �                      @        �       �                    �?$�q-�?	             *@        �       �                   `3@؇���X�?             @        ������������������������       �                     @        �       �                 03�7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        �       �                    @����E��?9            �V@       �       �                   �@@v�2t5�?5            �T@       �       �                 �|�=@҄��?)            �P@       �       �                     @�q�q��?             H@        ������������������������       �        	             .@        �       �                    @�q�q�?            �@@        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���7@����X�?             <@       �       �                    @r�q��?             2@        ������������������������       �                     @        �       �                    5@d}h���?	             ,@        �       �                  S%/@      �?             @        ������������������������       �                     �?        �       �                    +@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �/@ףp=
�?             $@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @      �?             $@        ������������������������       �                     @        �       �                 ��T?@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @D@�q�q�?             2@       �       �                    �?      �?	             0@        �       �                   �>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                      @        �       �                     @     ��?             0@       �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        �       �                    *@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @C@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �                          �?      �?J             ]@                                 !@@	tbA@�?)            @Q@        ������������������������       �                     �?        ������������������������       �        (             Q@              $                  @I@��C���?!            �G@                             `�>P@�Q����?             D@              
                �!fK@"pc�
�?             &@                              `�iJ@���Q��?             @        ������������������������       �                      @              	                   @@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @              #                p�w@J�8���?             =@             "                    �?R�}e�.�?             :@             !                   �?�X����?             6@                                 �?      �?             4@                               @G@�t����?             1@                               �9@r�q��?	             (@        ������������������������       �                     @                              �w|c@      �?              @                                �?�q�q�?             @        ������������������������       �                     �?                              03�U@z�G�z�?             @        ������������������������       �                     @                                �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                 �?���Q��?             @                               �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �*       h�h))��}�(h,h/h0M%KK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?R���Q�?���Q��?�?<<<<<<�?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�N���K�?]Ų����?��:m��?0��b�/�?�q�q�?r�q��?y�5���?Cy�5��?�������?ZZZZZZ�?              �?�؉�؉�?ى�؉��?F]t�E�?/�袋.�?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?              �?      �?              �?              �?      �?              �?      �?        UUUUUU�?�������?l�l��?��O��O�?�������?�������?              �?�?<<<<<<�?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?n۶m۶�?              �?      �?        ���Q��?R���Q�?              �?      �?      �?�������?UUUUUU�?�������?�������?      �?              �?      �?              �?      �?              �?        �������?�������?              �?�q�q�?�q�q�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �ҵ8f�?�iQR?δ?�q�q�?�q�q�?      �?        <<<<<<�?�?�������?UUUUUU�?�q�q�?�q�q�?;�;��?;�;��?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?        9��8���?�q�q�?�������?�?      �?              �?      �?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?        ��!:ܟ�?���.�?�؉�؉�?;�;��?�G�z�?���Q��?�Kh/��?h/�����?      �?        �k(���?(�����?333333�?�������?      �?      �?      �?        >����?|���?]t�E�?F]t�E�?      �?        <<<<<<�?�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?        ��Ǐ?�?����?�q�q�?�q�q�?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?             ��?      �?      �?        ��8��8�?�q�q�?      �?        �������?333333�?              �?��[��[�?�A�A�?F]t�E�?F]t�E�?�������?�?      �?      �?      �?                      �?      �?              �?        ------�?�������?UUUUUU�?UUUUUU�?�������?�������?      �?              �?      �?              �?�m۶m��?�$I�$I�?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?      �?        �a�a�?��y��y�?      �?        �������?�������?�$I�$I�?�m۶m��?              �?      �?              �?              �?        �0�0�?z��y���?O	� O�?b�־a�?333333�?�������?�������?ffffff�?      �?        �������?ZZZZZZ�?      �?      �?              �?vb'vb'�?;�;��?      �?      �?              �?�������?�������?      �?                      �?      �?              �?        颋.���?/�袋.�?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?                      �?h/�����?�Kh/��?              �?d!Y�B�?ӛ���7�?              �?�$I�$I�?�m۶m��?      �?                      �?�����?5�wL��?F]t�E�?t�E]t�?�a�a�?��y��y�?m��&�l�?'�l��&�?�؉�؉�?�;�;�?333333�?�������?              �?      �?      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?�������?333333�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?      �?        �������?�?      �?        �������?�?      �?        �؉�؉�?;�;��?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?                      �?      �?        }�'}�'�?�l�l�?�ڕ�]��?��+Q��?N6�d�M�?�d�M6��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?        �$I�$I�?�m۶m��?UUUUUU�?�������?              �?۶m۶m�?I�$I�$�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?�������?�������?      �?                      �?              �?      �?      �?              �?�������?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?      �?�q�q�?r�q��?              �?�������?�������?              �?      �?              �?              �?      �?              �?      �?              �?      �?ہ�v`��?�%~F��?      �?                      �?L� &W�?g���Q��?�������?ffffff�?F]t�E�?/�袋.�?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�rO#,��?|a���?'vb'vb�?�;�;�?�E]t��?]t�E]�?      �?      �?�������?�������?�������?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?              �?      �?              �?      �?              �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�-#hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                  x#J@ʡ�;S��?�           8�@              W                    �?V������?l           ��@               V                    @���i!��?l            `f@              7                    �?�q�q�?i            `e@                                  �?
�ۓQ{�?D            @\@                                X��C@ >�֕�?            �A@                                   @г�wY;�?             A@        ������������������������       �                      @        	       
                 �|Y8@ ��WV�?             :@        ������������������������       �                      @                                   �?�X�<ݺ?             2@        ������������������������       �                     �?                                 ��@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     �?                                  �#@�{ /h��?+            �S@                                  �5@���!pc�?             6@                                xF� @�q�q�?             @                                 �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                ���@      �?	             0@                                �|Y:@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �9@@4և���?             ,@       ������������������������       �                      @                                �?�@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        !       (                   �;@4և����?             L@        "       #                 pF%@�q�q�?	             8@        ������������������������       �                     (@        $       %                    7@r�q��?             (@        ������������������������       �                     @        &       '                   �7@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        )       4                     @     ��?             @@       *       -                 `f&'@ 	��p�?             =@        +       ,                   �J@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        .       /                   �E@�nkK�?             7@       ������������������������       �        	             0@        0       1                  ��9@؇���X�?             @       ������������������������       �                     @        2       3                   @H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        5       6                 ��1@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        8       E                    �?П[;U��?%             M@       9       :                     @b�2�tk�?             B@        ������������������������       �                     &@        ;       <                    @� �	��?             9@        ������������������������       �                     @        =       @                   �*@�z�G��?             4@        >       ?                    <@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        A       B                 `v�5@     ��?             0@        ������������������������       �                      @        C       D                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        F       I                    �?�eP*L��?             6@        G       H                 ��i<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        J       K                     @b�2�tk�?             2@        ������������������������       �                     @        L       O                    @8�Z$���?	             *@        M       N                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        P       Q                    ,@�C��2(�?             &@       ������������������������       �                     @        R       S                    �?      �?             @        ������������������������       �                      @        T       U                  `/@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        X       m                     �?d��K�T�?            �y@        Y       Z                 �|�<@�99lMt�?            �C@        ������������������������       �                     @        [       ^                    �?<ݚ)�?             B@        \       ]                 X�l@@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        _       l                  i?@�z�G��?             >@       `       k                   @=@      �?             2@       a       j                 `f�;@X�Cc�?	             ,@       b       c                   �B@�eP*L��?             &@        ������������������������       �                     @        d       e                 ��:@      �?              @        ������������������������       �                      @        f       g                   @G@�q�q�?             @        ������������������������       �                      @        h       i                   �K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             (@        n       �                 �?�@�n�Ƌ��?�            `w@        o       �                 �|�=@��a��?O            @^@       p       �                    �?㺦���?<            @W@        q       x                   �<@�>4և��?             <@        r       w                   �5@�8��8��?             (@        s       t                 �{@z�G�z�?             @        ������������������������       �                      @        u       v                   �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        y       �                    �?      �?             0@       z       {                 ���@�z�G��?             $@        ������������������������       �                     @        |       }                   @@և���X�?             @       ������������������������       ����Q��?             @        ~                        �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 �Y�@r�q��?             @        ������������������������       �                     �?        �       �                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �?$@��ɉ�?*            @P@       �       �                 ��@�7��?            �C@       �       �                     @г�wY;�?             A@        ������������������������       �                     @        �       �                  Md@ 7���B�?             ;@        ������������������������       �                     ,@        �       �                 ���@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        �       �                 �|Y8@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     :@        ������������������������       �                     <@        �       �                    �?Ԉ���a�?�            �o@        �       �                   �;@      �?	             2@       �       �                 �&2.@ףp=
�?             $@        �       �                 �&�)@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 @3�@H!s��?�            `m@        �       �                   �?@      �?             ,@       �       �                    :@����X�?             @       �       �                   �4@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �A@����X�?             @        ������������������������       �                      @        ������������������������       ����Q��?             @        �       �                    �?��[��?�            �k@       �       �                    �?t�G����?b            �e@        �       �                   `3@      �?             @        ������������������������       �                     �?        �       �                 03�7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     @ؙ/,T�?_             e@        �       �                   �*@     �?(             P@       �       �                   @A@$�q-�?            �C@       �       �                   @@@�����H�?             ;@       �       �                    &@$�q-�?             :@        �       �                    5@�����H�?             "@        ������������������������       �      �?             @        ������������������������       �                     @        �       �                   �(@�IєX�?             1@        ������������������������       �                     @        �       �                 �|�<@@4և���?
             ,@       ������������������������       �                     "@        �       �                 �|�=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             (@        ������������������������       �                     9@        �       �                 �|Y=@$�q-�?7             Z@       �       �                   �:@��� ��?             O@       �       �                   �3@      �?             H@        �       �                    2@��2(&�?             6@       �       �                 pf� @$�q-�?             *@        ������������������������       �z�G�z�?             @        ������������������������       �                      @        �       �                 `�8"@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     :@        �       �                 0S%"@X�Cc�?             ,@        �       �                 pf� @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���)@�<ݚ�?             "@       �       �                   �<@����X�?             @        ������������������������       �                     @        �       �                 ���"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     E@        �       �                 ��&@ \� ���?!            �H@        ������������������������       �                     @        �       �                    :@�3Ea�$�?              G@        �       �                    �?�LQ�1	�?             7@        ������������������������       �                     @        �       �                 03{3@���Q��?             4@        �       �                    0@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                 ���7@�	j*D�?	             *@       �       �                    �?�<ݚ�?             "@        ������������������������       �                     @        �       �                   �1@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                 ���A@�nkK�?             7@        ������������������������       �                     &@        �       �                   �C@�8��8��?             (@        �       �                   �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?�%~^��?K            �]@       �       �                  "�b@�Z��L��?+            �Q@       �       �                 ���Q@h㱪��?"            �K@        �       �                 @3[Q@؇���X�?             ,@       ������������������������       �        	             (@        ������������������������       �                      @        ������������������������       �                    �D@        �       �                    !@      �?	             0@        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �1@�q���?              H@        ������������������������       �                     @        �       �                   �8@�K��&�?            �E@        ������������������������       �                     @        �                          �?�\��N��?             C@       �       �                   �;@��}*_��?             ;@        ������������������������       �                     @                               `f^@�q�q�?             8@                               �H@      �?             4@                             `�iJ@      �?             0@        ������������������������       �                     �?                              �!fK@���Q��?             .@        ������������������������       �                     �?                              �|Y>@X�Cc�?
             ,@        ������������������������       �                     @              	                   �?"pc�
�?             &@        ������������������������       �                     @        
                           @���Q��?             @                             03�M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                 �?�C��2(�?             &@                             pU�t@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������N���I5�?d�~`l��?�g�`�|�?o0E>��?�D�H=�?�݇[@a�?UUUUUU�?UUUUUU�?��Ź��?2�s�8�?�A�A�?��+��+�?�?�?              �?;�;��?O��N���?              �?�q�q�?��8��8�?              �?�?�?      �?                      �?      �?        �|˷|��?�A�A�?F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?              �?      �?      �?      �?              �?      �?        n۶m۶�?�$I�$I�?      �?        �������?UUUUUU�?      �?                      �?n۶m۶�?%I�$I��?�������?�������?              �?�������?UUUUUU�?      �?        �m۶m��?�$I�$I�?      �?                      �?      �?      �?�{a���?������?UUUUUU�?�������?              �?      �?        d!Y�B�?�Mozӛ�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ��=���?�{a���?9��8���?�8��8��?              �?�Q����?)\���(�?              �?ffffff�?333333�?      �?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?        t�E]t�?]t�E�?      �?      �?      �?                      �?�8��8��?9��8���?              �?;�;��?;�;��?      �?      �?      �?                      �?]t�E�?F]t�E�?      �?              �?      �?      �?              �?      �?              �?      �?              �?        z��N52�?"�*7�?5H�4H��?�o��o��?              �?��8��8�?�8��8��?UUUUUU�?UUUUUU�?              �?      �?        ffffff�?333333�?      �?      �?%I�$I��?�m۶m��?t�E]t�?]t�E�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?      �?        ��X͞��?n�ʄm�?��2(&�?���|���?�]v�e��?EM4�D�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?333333�?�������?      �?      �?              �?      �?        �������?UUUUUU�?      �?        �������?�������?              �?      �?        ?�?��? �����?��[��[�?�A�A�?�?�?      �?        	�%����?h/�����?      �?        �؉�؉�?;�;��?              �?      �?        �������?�������?      �?              �?      �?      �?              �?        ���Sq��?�0�:��?      �?      �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        "c�]~��?ysB�n�?      �?      �?�$I�$I�?�m۶m��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�m۶m��?�$I�$I�?      �?        333333�?�������?�Ma�Ma�?�����?eMYS֔�?֔5eMY�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        z��y���?1�0ð?     ��?      �?�؉�؉�?;�;��?�q�q�?�q�q�?�؉�؉�?;�;��?�q�q�?�q�q�?      �?      �?      �?        �?�?      �?        n۶m۶�?�$I�$I�?      �?        �������?�������?              �?      �?                      �?      �?              �?        �؉�؉�?;�;��?�{����?�B!��?      �?      �?��.���?t�E]t�?�؉�؉�?;�;��?�������?�������?      �?        9��8���?�q�q�?              �?      �?              �?        %I�$I��?�m۶m��?�������?333333�?      �?                      �?9��8���?�q�q�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        
^N��)�?և���X�?              �?����7��?��,d!�?Nozӛ��?d!Y�B�?      �?        333333�?�������?۶m۶m�?�$I�$I�?              �?      �?        vb'vb'�?;�;��?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �Mozӛ�?d!Y�B�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        Rv�Qv��?�D �D �?��Vؼ?���.�d�?��)A��?־a���?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?      �?      �?                      �?�������?�������?              �?��)kʚ�?���)k��?      �?        y�5���?�5��P�?B{	�%��?_B{	�%�?              �?�������?�������?      �?      �?      �?      �?              �?�������?333333�?      �?        �m۶m��?%I�$I��?      �?        F]t�E�?/�袋.�?              �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ5�;5hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       f                     @�3)0�F�?�           8�@                                  �:@�G��l��?�            �s@                                   �?t���-��?:            �U@                                   �?H�z�G�?             D@        ������������������������       �                     1@                                   <@��+7��?             7@                                  5@�C��2(�?
             &@               	                   �2@r�q��?             @       ������������������������       �                     @        
                          �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?�q�q�?             (@                               �U�X@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                  �(@=QcG��?            �G@        ������������������������       �                      @                                ��f`@����?�?            �F@       ������������������������       �                     B@                                   !@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @               /                    �?~�І�^�?�            �l@                                  �;@�<p���?4            �T@                                   �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @               .                    �?`2U0*��?2            �R@               !                   �E@0G���ջ?%             J@       ������������������������       �                     A@        "       -                 ��A@r�q��?             2@        #       ,                 ���;@      �?              @       $       +                 `fF:@����X�?             @       %       &                   @F@���Q��?             @        ������������������������       �                     �?        '       *                    (@      �?             @       (       )                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     7@        0       ?                 ��D:@��-*�?_            @b@        1       >                   @A@�����?+            �P@       2       3                     �?�C��2(�?            �@@        ������������������������       �                     @        4       5                 �|Y=@ �Cc}�?             <@        ������������������������       �                     @        6       7                   �'@؇���X�?             5@        ������������������������       �                      @        8       =                 ��,@�θ�?
             *@        9       :                 �|�=@      �?             @        ������������������������       �                      @        ;       <                    @@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     A@        @       Q                    �?��It��?4            �S@        A       P                     �?д>��C�?             =@       B       O                 �UcV@���B���?             :@       C       N                    �?     ��?             0@       D       M                 @�6M@�n_Y�K�?	             *@       E       L                 p�i@@z�G�z�?             $@       F       K                    H@�q�q�?             @       G       H                 ��2>@�q�q�?             @        ������������������������       �                     �?        I       J                  �>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        R       e                     �?�w��#��?"             I@       S       X                 `f�;@r�qG�?              H@        T       U                    D@ףp=
�?             $@        ������������������������       �                     @        V       W                   @G@z�G�z�?             @        ������������������������       ��q�q�?             @        ������������������������       �                      @        Y       d                    �?���y4F�?             C@       Z       [                   �<@������?             A@        ������������������������       �                     @        \       c                   �Q@�חF�P�?             ?@       ]       b                 ���R@�r����?             >@       ^       _                   �H@ 7���B�?             ;@       ������������������������       �                     5@        `       a                   �J@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        g       �                    �?���!pc�?�            �x@        h       �                 03�:@vs�G��?I            �]@       i       |                    �?+Y���?E            @\@        j       o                 P��+@� ��1�?            �D@       k       l                    �?$�q-�?             :@        ������������������������       �                     @        m       n                    �?�����?             5@       ������������������������       �        
             3@        ������������������������       �                      @        p       s                    �?���Q��?
             .@        q       r                  S�-@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        t       u                 03�-@      �?              @        ������������������������       �                     @        v       w                    �?      �?             @        ������������������������       �                     �?        x       {                    @�q�q�?             @       y       z                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        }       �                    �?�E��ӭ�?-             R@       ~       �                    �?�G�z��?             D@              �                 �|Y=@h+�v:�?             A@        �       �                 �&�)@��Q��?
             4@       �       �                 ���@؇���X�?             ,@        �       �                   �7@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �5@�C��2(�?             &@        ������������������������       �                     @        �       �                   @@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �0@r�q��?             @        ������������������������       �                     @        �       �                   �2@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                   �2@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @@       �       �                 X��A@`Jj��?             ?@       �       �                 ���@�>����?             ;@        ������������������������       �                     "@        �       �                   @'@�����H�?             2@       ������������������������       �"pc�
�?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��PBKP�?�            `q@        �       �                    �?�s��:��?3             S@       �       �                    @��k��?!            �J@        ������������������������       �                     @        �       �                    *@      �?             H@        �       �                    @r�q��?             @       �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 03�1@��6���?             E@       �       �                   �D@b�2�tk�?             B@       �       �                  �#@ҳ�wY;�?             A@       �       �                   �@�G��l��?             5@        �       �                 �|Y:@�	j*D�?             *@       �       �                 pf�@"pc�
�?             &@        ������������������������       �                     @        �       �                 �&B@�q�q�?             @       �       �                    4@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �*@8�Z$���?	             *@        ������������������������       �                     @        �       �                 �|�<@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 `fV6@r�q��?             @        �       �                   �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @��<b���?             7@       �       �                    @�GN�z�?             6@        �       �                    @      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �6@      �?             0@        ������������������������       �                      @        �       �                 ��p@@      �?              @        �       �                   @C@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       
                   �?8Fb����?�            @i@       �                       �T)D@��0��?m            �e@       �                         �C@���Cu��?j            �d@       �       �                 �|�=@����1�?`            @b@       �       �                 pf� @,Z0R�?J             ]@       �       �                   �0@$��$�L�?6            �S@        ������������������������       �                     �?        �       �                 ��) @�:�^���?5            �S@       �       �                   �8@`-�I�w�?4             S@        �       �                   �7@��-�=��?            �C@       �       �                 @3�@�IєX�?             A@       �       �                   �3@Pa�	�?            �@@        ������������������������       �        	             0@        �       �                 �?�@�IєX�?             1@       ������������������������       �        
             ,@        �       �                   �4@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 03@���Q��?             @       �       �                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                 �?$@�?�|�?            �B@        �       �                 pf�@�����H�?             "@       ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     <@        ������������������������       �                      @        �       �                 ���#@�?�|�?            �B@       �       �                 ���"@���7�?             6@       ������������������������       �                     *@        �       �                   �<@�����H�?             "@        ������������������������       �                     @        �       �                 �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             .@        �       �                   @@@r�q��?             >@        �       �                 �?�@�	j*D�?	             *@        ������������������������       �                     @        �       �                 ��Y)@���Q��?             $@       �       �                 �̌!@      �?              @       �       �                 @3�@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @                                 @C@�IєX�?             1@       ������������������������       �        
             ,@                              ��	0@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �        
             5@              	                �|�>@���Q��?             @                             �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                 @�r����?             >@                              @3�4@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     2@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������Rl���?�[�'��?��y��y�?1�0��?��֡�l�?�L�Ȥ�?333333�?ffffff�?              �?zӛ����?Y�B��?]t�E�?F]t�E�?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?        �������?�������?�$I�$I�?�m۶m��?              �?      �?              �?        AL� &W�?x6�;��?      �?        l�l��?��I��I�?              �?�q�q�?�q�q�?      �?                      �?�#���>�?$���>��?�����?}���|�?۶m۶m�?�$I�$I�?              �?      �?        {�G�z�?���Q��?�؉�؉�?vb'vb'�?              �?UUUUUU�?�������?      �?      �?�$I�$I�?�m۶m��?�������?333333�?      �?              �?      �?      �?      �?              �?      �?                      �?              �?      �?                      �?              �?T�P�B��?�^�z���?g��1��?���@��?]t�E�?F]t�E�?      �?        %I�$I��?۶m۶m�?      �?        ۶m۶m�?�$I�$I�?      �?        ى�؉��?�؉�؉�?      �?      �?              �?      �?      �?      �?              �?      �?      �?              �?        -n����?�#{���?a���{�?|a���?��؉���?ى�؉��?      �?      �?;�;��?ى�؉��?�������?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?                      �?      �?              �?              �?        ��Q��?��(\���?�������?�������?�������?�������?              �?�������?�������?UUUUUU�?UUUUUU�?              �?6��P^C�?(������?xxxxxx�?�?              �?�Zk����?��RJ)��?�������?�?	�%����?h/�����?      �?        �������?UUUUUU�?              �?      �?                      �?              �?      �?              �?        F]t�E�?t�E]t�?���؊��?�N��?��	���?H���?������?������?;�;��?�؉�؉�?              �?�a�a�?=��<���?              �?      �?        �������?333333�?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?�q�q�?r�q��?�������?�������?�������?xxxxxx�?ffffff�?�������?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?]t�E�?              �?      �?      �?      �?                      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?      �?                      �?      �?      �?���{��?�B!��?�Kh/��?h/�����?      �?        �q�q�?�q�q�?/�袋.�?F]t�E�?      �?              �?              �?              �?        �n��G��?�Eΰ�R�?��k(��?�k(���?"5�x+��?oe�Cj��?              �?      �?      �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        =��<���?b�a��?9��8���?�8��8��?�������?�������?��y��y�?1�0��?;�;��?vb'vb'�?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?              �?      �?      �?                      �?;�;��?;�;��?              �?      �?      �?      �?                      �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��,d!�?��Moz��?�袋.��?]t�E�?      �?      �?      �?                      �?      �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        =�]?[��?�&��?6eMYS��?S֔5eM�?�8��>Q�?@:�2	v�?�Ν;w��?Ĉ#F��?�FX�i��?	�=��ܳ?��]-n��?�3���?              �?� � �?�o��o��?Q^Cy��?y�5�װ?}˷|˷�?�A�A�?�?�?|���?|���?      �?        �?�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        *�Y7�"�?к����?�q�q�?�q�q�?      �?              �?      �?      �?                      �?*�Y7�"�?к����?�.�袋�?F]t�E�?      �?        �q�q�?�q�q�?      �?        �������?�������?              �?      �?              �?        �������?UUUUUU�?vb'vb'�?;�;��?      �?        333333�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �?�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�?UUUUUU�?UUUUUU�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJi4�hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       f                    �?H���I�?�           8�@               e                    @��j!D��?�            `n@              &                    �?�aʬ��?�            �m@                                   �?ףp=
�?8             T@                                   @�NW���?(            �J@                                  �?h�����?             <@              
                     �? ��WV�?             :@              	                 03�=@ �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                      @        ������������������������       �                      @                                  �-@H%u��?             9@                                  �,@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                �|�9@���}<S�?             7@        ������������������������       �                     @                                   �?�����H�?             2@                                ��%@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                ���@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �        
             ,@                                   @PN��T'�?             ;@        ������������������������       �                     @                                    @z�G�z�?             4@       ������������������������       �                     ,@               %                    @�q�q�?             @                                �|�7@z�G�z�?             @        ������������������������       �                      @        !       $                    �?�q�q�?             @       "       #                 X��B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        '       <                 Ь�#@"��5��?f            �c@        (       /                   �@�n_Y�K�?             :@        )       .                 �|�;@�q�q�?             "@       *       +                 ���@؇���X�?             @        ������������������������       �                     @        ,       -                    4@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        0       1                 �?�@������?
             1@        ������������������������       �                     @        2       3                    3@����X�?	             ,@        ������������������������       �                      @        4       ;                 `��!@r�q��?             (@       5       :                 �|Y>@      �?              @       6       9                 @3�@؇���X�?             @       7       8                   �8@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        =       R                     @���4Z��?T            ``@       >       A                    @��r
'��?:            @W@        ?       @                     �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        B       C                     �?�:�^���?8            �V@        ������������������������       �                     @@        D       Q                    �?\-��p�?"             M@       E       F                 `f�)@r٣����?            �@@        ������������������������       �                     $@        G       N                   �E@�LQ�1	�?             7@       H       M                   �7@�<ݚ�?             2@       I       J                   �;@���Q��?	             $@        ������������������������       �                     @        K       L                   �B@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        O       P                   @F@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     9@        S       `                 03�1@p�ݯ��?             C@        T       Y                   �*@�E��ӭ�?             2@        U       X                 ��&@      �?              @        V       W                    4@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        Z       [                 ��Y.@���Q��?             $@        ������������������������       �                     @        \       _                    �?؇���X�?             @       ]       ^                 �|�;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        a       d                  �7@P���Q�?             4@        b       c                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             *@        ������������������������       �                     @        g       �                 ��i=@�Ն���?(           @}@       h       �                    �?�&�TA�?�             w@        i       �                    �?�θ�?/            �S@       j       {                 ��i @�D��?            �H@       k       l                 03S@��G���?            �B@        ������������������������       �                     @        m       x                   @@H�V�e��?             A@       n       q                 ���@      �?             8@        o       p                 �|�9@      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        r       s                   @8@      �?             (@        ������������������������       �                      @        t       u                 �|=@ףp=
�?             $@        ������������������������       �                     �?        v       w                 �|�=@�����H�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        y       z                 �|Y=@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        |       �                  A7@      �?	             (@       }       ~                     @�q�q�?             "@        ������������������������       �                      @               �                 �|Y?@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ;@д>��C�?             =@        ������������������������       �                     $@        �       �                     @�d�����?             3@        ������������������������       �                     �?        �       �                 �|Y=@�E��ӭ�?             2@        ������������������������       �                      @        �       �                   `3@     ��?             0@       �       �                   @'@�r����?             .@       �       �                 �Y�@"pc�
�?             &@        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 `ff:@DK{22�?�             r@       �       �                     �?�Km�a̾?�            �q@        ������������������������       �                     @        �       �                    �?`�BX�l�?�             q@       �       �                     @,(��?�            �o@        �       �                 `f�)@$Q�q�?'            �O@        ������������������������       �                     7@        �       �                 �|Y=@ףp=
�?             D@        ������������������������       �                     *@        �       �                 �|�=@PN��T'�?             ;@        ������������������������       �                     �?        �       �                   �*@ȵHPS!�?             :@       �       �                    @@     ��?	             0@        ������������������������       �                     @        �       �                   @B@�z�G��?             $@        ������������������������       ��q�q�?             @        �       �                   �F@؇���X�?             @       �       �                   @D@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     $@        �       �                 ���!@�F�l���?w            �g@       �       �                 ��) @��F��?`            `c@       �       �                   �2@�t:ɨ�?S            �`@        �       �                 ���@z�G�z�?             $@       ������������������������       �                     @        �       �                    1@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                 �?$@ ;=֦��?L            �^@        �       �                 �|�?@�}�+r��?             C@       �       �                 ���@HP�s��?             9@       �       �                    7@���N8�?             5@        ������������������������       �                      @        �       �                   �8@$�q-�?             *@        �       �                 �&b@؇���X�?             @        ������������������������       �                     @        �       �                 `fF@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|Y8@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �        
             *@        �       �                 @3�@ ��N8�?1             U@       �       �                   �B@`Ql�R�?            �G@       ������������������������       �                     E@        �       �                 �?�@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                    �B@        �       �                   �:@�LQ�1	�?             7@       ������������������������       �                     *@        �       �                 �|Y<@�z�G��?             $@        ������������������������       �                      @        �       �                 pF� @      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     B@        �       �                    �?�z�G��?             4@       �       �                    (@�E��ӭ�?             2@       �       �                    @X�<ݚ�?             "@        �       �                 ף�?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                   �4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 `f�;@�z�G��?             $@       �       �                 �|�<@�q�q�?             "@        ������������������������       �                     �?        �       �                 �|�?@      �?              @        ������������������������       �                      @        �       �                   �C@�q�q�?             @        ������������������������       �                     �?        �       �                    H@z�G�z�?             @        ������������������������       �                      @        �       �                   �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 03#?@�w��#��?A             Y@        �       �                    �?      �?
             0@       �       �                  I>@؇���X�?	             ,@       �       �                    �?�q�q�?             @       �       �                     �?�q�q�?             @       �       �                 X��E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    @0,Tg��?7             U@        �       �                     @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          �?�6i����?3            �S@       �                          �?�q����?#            �J@        �       �                 м�J@�q�q�?	             (@        ������������������������       �                      @        �                          �H@      �?             $@       �       �                 X�,@@����X�?             @        �       �                 0�HU@�q�q�?             @        ������������������������       �                     �?        �       �                 Ȫ�c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  @���� �?            �D@                             ���[@��hJ,�?             A@                                �?��a�n`�?             ?@        ������������������������       �                     �?              	                  �<@ףp=
�?             >@                              `f�D@      �?              @        ������������������������       �                      @        ������������������������       �                     @        
                         A@���7�?             6@                              �|Y>@�C��2(�?             &@        ������������������������       �                     @                                @K@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             &@                               �6f@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 ;@؇���X�?             @        ������������������������       �                     @                                 >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 �?$�q-�?             :@                                �7@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     1@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������Q�Ȟ���?^-n����?�F�� ��?�\��o��?��sI,S�?��4+�?�������?�������?�x+�R�?萚`���?�$I�$I�?�m۶m��?;�;��?O��N���?UUUUUU�?�������?      �?                      �?              �?              �?���Q��?)\���(�?      �?      �?              �?      �?        d!Y�B�?ӛ���7�?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?        �?�������?      �?                      �?h/�����?&���^B�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?����a�?�:�2��?;�;��?ى�؉��?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        xxxxxx�?�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?      �?        Ls�U��?ZF�ձ�?�n�ᆻ?�<��#��?UUUUUU�?UUUUUU�?      �?                      �?l�l��?}�'}�'�?              �?�{a���?a����?|���?>���>�?              �?d!Y�B�?Nozӛ��?�q�q�?9��8���?�������?333333�?      �?        �$I�$I�?۶m۶m�?              �?      �?                      �?�������?�������?      �?                      �?              �?^Cy�5�?Cy�5��?r�q��?�q�q�?      �?      �?      �?      �?              �?      �?                      �?�������?333333�?      �?        �$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?ffffff�?�������?۶m۶m�?�$I�$I�?      �?                      �?      �?              �?        #0#0�?t?�s?��?�Mozӛ�?���,d!�?ى�؉��?�؉�؉�?������??4և���?#�u�)��?v�)�Y7�?      �?        iiiiii�?ZZZZZZ�?      �?      �?      �?      �?              �?      �?              �?      �?              �?�������?�������?      �?        �q�q�?�q�q�?      �?      �?      �?        �������?�������?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?        a���{�?|a���?      �?        Cy�5��?y�5���?      �?        �q�q�?r�q��?              �?      �?      �?�������?�?/�袋.�?F]t�E�?      �?              �?      �?      �?                      �?���Dɮ�?^�(ٵ��?_�_��?PuPu�?      �?        �������?��;�HѰ?�����|�?��`0�?~��}���?AA�?      �?        �������?�������?      �?        &���^B�?h/�����?              �?��N��N�?�؉�؉�?      �?      �?      �?        ffffff�?333333�?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?        L�:,��?:kP<�q�?Y���/Y�?mЦm�?�&�l���?e�M6�d�?�������?�������?      �?              �?      �?UUUUUU�?UUUUUU�?              �?�%C��6�?XG��).�?�5��P�?(�����?q=
ףp�?{�G�z�?��y��y�?�a�a�?      �?        �؉�؉�?;�;��?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?              �?      �?      �?        �y��y��?�a�a�?}g���Q�?W�+�ɕ?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?      �?        ��Moz��?Y�B��?      �?        ffffff�?333333�?              �?      �?      �?              �?      �?              �?        ffffff�?333333�?�q�q�?r�q��?�q�q�?r�q��?�������?�������?              �?      �?                      �?      �?              �?      �?              �?      �?        ffffff�?333333�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ��Q��?��(\���?      �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?              �?      �?        �y��y��?1�0��?�������?�������?              �?      �?        kq�w��?T:�g *�?�Cj��V�?�x+�R�?�������?�������?      �?              �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        jW�v%j�?,Q��+�?KKKKKK�?�������?�s�9��?�c�1Ƹ?      �?        �������?�������?      �?      �?              �?      �?        �.�袋�?F]t�E�?]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?�؉�؉�?;�;��?9��8���?�q�q�?              �?      �?              �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ThG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       �                   �R@<C�`��?�           8�@              Y                    �?8	C)��?�           ��@               V                 pfP@2X��ʑ�?o            �e@              C                 Ь�9@������?k            �d@                                   @3k���?L            @\@                                   �?�ݜ�?            �C@        ������������������������       �                      @                                  �+@�חF�P�?             ?@       	                          �'@���y4F�?             3@        
                          �J@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?                                   ;@�q�q�?             "@        ������������������������       �                      @                                   B@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  @4@�8��8��?	             (@        ������������������������       �                     @                                   �?z�G�z�?             @                                   ?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                    '@��%��?4            �R@                                   �?�z�G��?             $@                                  �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   @؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        !       B                  ��8@     8�?.             P@       "       #                   �3@�0u��A�?,             N@        ������������������������       �                      @        $       9                 ��.@��WV��?%             J@       %       ,                 �|�<@�s��:��?             C@        &       '                 ��@ҳ�wY;�?             1@        ������������������������       �                     @        (       )                    �?�8��8��?             (@       ������������������������       �                     "@        *       +                   �*@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        -       8                    �?�G��l��?             5@       .       /                 ���@ҳ�wY;�?             1@        ������������������������       �                      @        0       7                 ���*@������?             .@       1       6                    C@8�Z$���?             *@       2       3                  ��@�8��8��?
             (@       ������������������������       �                     "@        4       5                 ��� @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        :       ;                 �|�=@؇���X�?
             ,@       ������������������������       �                     $@        <       =                   �>@      �?             @        ������������������������       �                     �?        >       ?                 ���0@�q�q�?             @        ������������������������       �                     �?        @       A                 03C3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        D       Q                    @@�0�!��?            �I@       E       L                    '@�:�^���?            �F@        F       K                    !@�z�G��?             $@       G       H                    @      �?              @        ������������������������       �                     @        I       J                     @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        M       N                 03;<@��?^�k�?            �A@        ������������������������       �        	             3@        O       P                 0Cd=@      �?
             0@        ������������������������       �                     �?        ������������������������       �        	             .@        R       U                 ��p@@r�q��?             @        S       T                   @C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        W       X                 X�l@@      �?              @       ������������������������       �                     @        ������������������������       �                      @        Z       �                 �?�@���6�.�?           �|@        [       �                    �?���g�X�?X            `b@       \       k                   �8@ )�y���?W             b@        ]       d                    �?؇���X�?            �A@        ^       a                    5@      �?              @        _       `                 �{@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        b       c                 ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        e       j                 ���@�>����?             ;@        f       g                    7@����X�?             @        ������������������������       �                     @        h       i                 �&b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     4@        l       u                    �?Ц�f*�?B            �[@        m       n                 �|=@P���Q�?             4@        ������������������������       �                     @        o       t                 �|�=@$�q-�?	             *@       p       q                 ���@�����H�?             "@        ������������������������       �                     @        r       s                   @@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        ������������������������       �                     @        v       w                    �?����?�?7            �V@        ������������������������       �                     5@        x       y                    ?@��.N"Ҭ?*            @Q@       ������������������������       �                    �D@        z       {                 �&B@@4և���?             <@       ������������������������       �                     6@        |                           A@�q�q�?             @        }       ~                   �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 @3�@�4 )��?�            ps@        �       �                   �4@��
ц��?	             *@        ������������������������       �      �?             @        �       �                   �=@�q�q�?             "@        ������������������������       �                     @        �       �                   �?@���Q��?             @        ������������������������       �                     �?        �       �                   �A@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                    �?u�����?�            �r@       �       �                 `fF:@�Q��k�?�             n@       �       �                    �?$�Q�\�?j             e@        �       �                     @���!pc�?	             &@        ������������������������       �                      @        �       �                   �:@�q�q�?             "@        �       �                 �y.@      �?             @        ������������������������       �                     �?        �       �                   �2@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                     @�d	���?a            �c@        �       �                   �*@ �h�7W�?"            �J@       �       �                 `f�)@     ��?             @@       �       �                   �7@���N8�?             5@        �       �                    &@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             0@        �       �                 �|�<@"pc�
�?	             &@       ������������������������       �                     @        �       �                 �|�=@���Q��?             @        ������������������������       �                     �?        �       �                    B@      �?             @        ������������������������       �                      @        �       �                    G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        �       �                 ���!@(N:!���??            @Z@       �       �                 @Q!@��x_F-�?             �I@       �       �                   �3@�T|n�q�?            �E@        �       �                 0S5 @      �?             (@       �       �                    1@���Q��?             $@        ������������������������       ����Q��?             @        �       �                   �2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                      @        �       �                 �|�=@�g�y��?             ?@       �       �                 ��) @P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                 �|Y<@      �?              @        �       �                    8@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �<@ 7���B�?             K@        ������������������������       �                     8@        �       �                    �?��S�ۿ?             >@        �       �                   `3@�C��2(�?             &@       ������������������������       �                     @        �       �                 03�7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 �|Y=@�}�+r��?             3@        �       �                 ���"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             1@        �       �                   �<@����O��?/            �Q@        �       �                    7@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?d��0u��?)             N@        �       �                   �@@������?             .@        ������������������������       �                     @        �       �                   @J@      �?              @       �       �                   �A@z�G�z�?             @        ������������������������       �                     @        �       �                  xCH@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                      @z�G�z�?            �F@       �       �                   �G@"pc�
�?             F@       �       �                 �|Y>@��a�n`�?             ?@        ������������������������       �                     &@        �       �                   �A@R���Q�?             4@        �       �                   @@@���Q��?             @       �       �                   @K@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �F@��S�ۿ?	             .@        �       �                 03�C@r�q��?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     "@        �       �                   �J@�n_Y�K�?             *@        �       �                   @I@����X�?             @        �       �                   �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�BbΊ�?#             M@        �       �                 X��@@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                    @��[�p�?            �G@        �       �                   �;@�q�q�?             .@       ������������������������       �                     "@        �       �                    �?r�q��?             @        �       �                 ��yE@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @@        �                          �?�Zl�i��?/            @T@       �                          �?Du9iH��?            �E@       �                           �?������?            �D@       ������������������������       �                    �@@                                 �?      �?              @                               �5@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                              hfzg@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        	      
                   �?�?�'�@�?             C@       ������������������������       �                     <@                                 �?      �?             $@                             ���[@      �?              @                               �D@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                               �6f@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub�������������܍�W�?/�F�JP�?�h��h��?S.�R.��?}A_��?}A_���?��+Q��?�v%jW��?zja���?�JO-���?�i�i�?\��[���?              �?��RJ)��?�Zk����?(������?6��P^C�?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?      �?                      �?              �?}���g�?���L�?ffffff�?333333�?UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?     ��?�������?�������?              �?��N��N�?��؉���?��k(��?�k(���?�������?�������?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��y��y�?1�0��?�������?�������?      �?        �?wwwwww�?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        �������?ZZZZZZ�?l�l��?}�'}�'�?333333�?ffffff�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �A�A�?_�_��?              �?      �?      �?      �?                      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?Ct�?�?���.�?��fG-B�?���+ݫ?q��<�?����?�?۶m۶m�?�$I�$I�?      �?      �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �Kh/��?h/�����?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        !O	� �?�־a�?ffffff�?�������?      �?        �؉�؉�?;�;��?�q�q�?�q�q�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?        ��I��I�?l�l��?      �?        �3J���?ہ�v`��?      �?        n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �C��?���̱�?�;�;�?�؉�؉�?      �?      �?UUUUUU�?UUUUUU�?      �?        �������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?!��*�3�?}0T�1�?�������?�������?)ݾ�z��?�	j*D�?F]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��JG��?�0���M�?��sHM0�?"5�x+��?      �?      �?��y��y�?�a�a�?�������?�������?              �?      �?              �?        /�袋.�?F]t�E�?      �?        333333�?�������?              �?      �?      �?      �?              �?      �?              �?      �?              �?        |�W|�W�?�A�A�?�������?�?���)k��?6eMYS��?      �?      �?�������?333333�?333333�?�������?�������?�������?              �?      �?      �?      �?        ��{���?�B!��?ffffff�?�������?      �?                      �?      �?              �?      �?�������?333333�?      �?                      �?      �?        	�%����?h/�����?      �?        �������?�?]t�E�?F]t�E�?      �?              �?      �?              �?      �?        �5��P�?(�����?      �?      �?      �?                      �?      �?         �
���?�]�����?t�E]t�?F]t�E�?      �?                      �?�?�������?wwwwww�?�?      �?              �?      �?�������?�������?              �?      �?      �?      �?                      �?      �?        �������?�������?/�袋.�?F]t�E�?�s�9��?�c�1Ƹ?      �?        333333�?333333�?333333�?�������?      �?      �?      �?                      �?              �?�������?�?�������?UUUUUU�?      �?      �?      �?              �?        ;�;��?ى�؉��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�{a��?���=��?t�E]t�?]t�E�?              �?      �?        �
br1�?m�w6�;�?UUUUUU�?UUUUUU�?              �?�������?UUUUUU�?      �?      �?              �?      �?              �?              �?        �����H�?�"e����?w�qGܱ?qG�w��?������?p>�cp�?              �?      �?      �?�$I�$I�?�m۶m��?      �?                      �?              �?      �?      �?      �?                      �?y�5���?������?              �?      �?      �?      �?      �?�������?�������?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ5�R/hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       8                    �?t�C�#��?�           8�@                                   �?T�7�s��?p            `e@                                   @ �\���?/            �S@                                  &@ ��WV�?.            �S@                                   @����X�?             @       ������������������������       �                     @        ������������������������       �                      @               	                 �|Y=@ ��PUp�?+            �Q@        ������������������������       �                     <@        
                        �|�=@ qP��B�?            �E@                                ���@P���Q�?             4@        ������������������������       �                     �?        ������������������������       �        
             3@        ������������������������       �                     7@        ������������������������       �                     �?               7                 �̾w@�W��?A             W@                               03s@
�GN��??             V@        ������������������������       �                     <@               6                    �?��0u���?)             N@              5                 p"�X@�BbΊ�?'             M@              4                    �?�t����?"            �I@              /                    �?      �?             D@                                  2@X�Cc�?             <@        ������������������������       �                      @               "                 �|Y=@�	j*D�?             :@               !                   �:@�eP*L��?             &@                               �0@�q�q�?             "@        ������������������������       �                     @                                Ȉ�P@���Q��?             @        ������������������������       �                      @                                   �8@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        #       $                    A@z�G�z�?             .@        ������������������������       �                     @        %       .                 ��O@      �?              @       &       -                   �A@����X�?             @       '       ,                     �?���Q��?             @       (       )                    <@      �?             @        ������������������������       �                     �?        *       +                 ��Y>@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        0       3                     @�q�q�?             (@       1       2                 ��UO@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        9       �                    �?<ݚ)�?N           ��@        :                           �?N§�r��?l            �f@       ;       Z                     @����&�?V            �`@       <       W                    L@���}<S�?7             W@       =       >                     �? 	��p�?4            �U@        ������������������������       �                     A@        ?       V                    �?���C��?!            �J@       @       K                   �2@�MI8d�?            �B@       A       B                    :@�C��2(�?             6@        ������������������������       �                     �?        C       J                   �*@���N8�?             5@       D       E                 `f�)@��S�ۿ?
             .@        ������������������������       �                     @        F       G                   �B@ףp=
�?             $@       ������������������������       �                      @        H       I                    D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        L       O                    <@������?	             .@        M       N                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        P       Q                   �7@�C��2(�?             &@        ������������������������       �                     �?        R       U                   �=@ףp=
�?             $@       S       T                   �E@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             0@        X       Y                     �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        [       `                    @�+��<��?            �E@        \       ]                    @      �?              @        ������������������������       �                     @        ^       _                 @3�2@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        a       b                 ���@^������?            �A@        ������������������������       �                      @        c       d                   �5@:ɨ��?            �@@        ������������������������       �                     @        e       p                 ��&@�n_Y�K�?             :@       f       o                    �?d}h���?             ,@       g       n                 03�!@      �?             (@       h       i                    8@�q�q�?             "@        ������������������������       �                      @        j       k                 �?�@؇���X�?             @       ������������������������       �                     @        l       m                   �9@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        q       z                    �?�q�q�?	             (@       r       y                 03�1@      �?             @       s       t                 @3�/@      �?             @        ������������������������       �                     �?        u       x                   �0@�q�q�?             @       v       w                 �|�;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        {       |                   �;@�q�q�?             @        ������������������������       �                     @        }       ~                 �|Y>@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                     @�L�lRT�?            �F@        �       �                 ���[@�8��8��?             (@       ������������������������       �                     "@        �       �                 ���i@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 `f�8@6YE�t�?            �@@        ������������������������       �                     @        �       �                    @��S�ۿ?             >@       ������������������������       �        
             8@        �       �                    @�q�q�?             @       �       �                 ��T?@      �?             @        ������������������������       �                     �?        �       �                 ���A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?<�Z��?�            �v@       �       �                 ��$:@ ��om��?�            ps@       �       �                 �?�@��Y�h9�?�            @o@        �       �                 ��@�O4R���?=            �Z@        ������������������������       �                    �I@        �       �                 �?$@h㱪��?            �K@        �       �                 �|�;@z�G�z�?             $@       ������������������������       �                     @        �       �                 X��I@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �F@        �       �                 @3�@8��8���?Z             b@        �       �                   �9@      �?             @        ������������������������       �                     �?        �       �                   �?@���Q��?             @        ������������������������       �                     �?        �       �                   �A@      �?             @       ������������������������       ��q�q�?             @        ������������������������       �                     �?        �       �                     @���}<S�?T            @a@        �       �                   �@@      �?"             H@       ������������������������       �                     =@        �       �                   @A@�S����?             3@        �       �                   �3@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        �       �                 �|Y=@ףp=
�?2            �V@       �       �                   �9@�������?             F@       �       �                 0S5 @؇���X�?            �A@        �       �                   �3@�q�q�?             (@        �       �                   �1@r�q��?             @       ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     7@        �       �                   �;@X�<ݚ�?             "@        ������������������������       �                      @        �       �                   �<@����X�?             @       ������������������������       �                     @        �       �                 �̌!@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     G@        �       �                     �?�'N��?)            �N@       �       �                  i?@"Ae���?#            �G@        �       �                    K@D�n�3�?             3@       �       �                   �<@      �?
             (@        ������������������������       �                     @        �       �                   @>@�q�q�?             "@       �       �                   �?@և���X�?             @        ������������������������       �                      @        �       �                    D@z�G�z�?             @        ������������������������       �                      @        �       �                   @G@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 `fF<@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 03�U@�>4և��?             <@       �       �                   @K@�LQ�1	�?             7@       �       �                 �|�<@z�G�z�?             .@        �       �                    7@      �?             @        ������������������������       �                     �?        �       �                 `f�D@�q�q�?             @        ������������������������       �                     �?        �       �                   �;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 0�J@�C��2(�?	             &@       ������������������������       �                     "@        �       �                 `�iJ@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                 X��@@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    ;@@4և���?             ,@        �       �                 ��?P@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 �̌4@ \� ���?"            �H@        �       �                 ���"@��
ц��?
             *@        ������������������������       �                     @        �       �                   �3@���Q��?	             $@       �       �                 ��L.@����X�?             @       �       �                    -@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                     @r�q��?             B@        �       �                 `��S@     ��?             0@       �       �                    �?"pc�
�?             &@       �       �                    :@����X�?             @        ������������������������       �                     �?        �       �                    0@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    5@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �                       ���A@P���Q�?             4@                               ��T?@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub��������������td�@�?��7a~�?�}��?p�}��?�3���?���7a�?;�;��?O��N���?�$I�$I�?�m۶m��?              �?      �?        ��V،?��ۥ���?              �?�}A_З?��}A�?�������?ffffff�?      �?                      �?              �?      �?        Y�B��?ӛ���7�?�E]t��?�袋.��?      �?        �������?""""""�?�{a��?���=��?�������?�������?      �?      �?%I�$I��?�m۶m��?              �?vb'vb'�?;�;��?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?              �?      �?�m۶m��?�$I�$I�?333333�?�������?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?�������?�������?9��8���?�q�q�?      �?                      �?              �?      �?              �?                      �?              �?��8��8�?�8��8��?[�[��?}�'}�'�?t��:W�?���M1j�?d!Y�B�?ӛ���7�?�{a���?������?              �?"5�x+��?\�琚`�?L�Ϻ��?��L���?F]t�E�?]t�E�?      �?        �a�a�?��y��y�?�?�������?              �?�������?�������?              �?      �?      �?      �?                      �?              �?�?wwwwww�?      �?      �?      �?                      �?F]t�E�?]t�E�?              �?�������?�������?�q�q�?�q�q�?              �?      �?                      �?              �?�������?333333�?              �?      �?        w�qG��?w�qG�?      �?      �?              �?      �?      �?              �?      �?        uPuP�?_�_��?              �?N6�d�M�?e�M6�d�?      �?        ;�;��?ى�؉��?I�$I�$�?۶m۶m�?      �?      �?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�I��I��?l�l��?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?'�l��&�?e�M6�d�?              �?�������?�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �>�>��?�[�[�?�]i��?�����?m������?�� �rh�?:�&oe�?�x+�R�?      �?        ־a���?��)A��?�������?�������?      �?              �?      �?              �?      �?              �?        �������?�������?      �?      �?      �?        �������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?ӛ���7�?d!Y�B�?      �?      �?      �?        (������?^Cy�5�?      �?      �?              �?      �?              �?        �������?�������?t�E]t�?/�袋.�?۶m۶m�?�$I�$I�?�������?�������?UUUUUU�?�������?      �?      �?              �?      �?              �?        r�q��?�q�q�?              �?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?      �?        �����?ާ�d��?�w6�;�?W�+���?(������?l(�����?      �?      �?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?              �?              �?�m۶m��?�$I�$I�?      �?                      �?�$I�$I�?�m۶m��?��Moz��?Y�B��?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        ]t�E�?F]t�E�?      �?              �?      �?              �?      �?              �?        333333�?�������?      �?                      �?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?              �?      �?              �?        
^N��)�?և���X�?�;�;�?�؉�؉�?      �?        �������?333333�?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?      �?      �?/�袋.�?F]t�E�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?              �?      �?              �?        �������?333333�?              �?      �?        ffffff�?�������?      �?      �?      �?                      �?      �?        ��       ubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�%hG        hNhG        hNh>Kh@KhAh))��}�(h,h/h0K��h2h3h4hVh<�h=Kub�              �?�B       hJhZhGC       ���R�h^Kh_hbKh))��}�(h,h/h0K��h2h3h4hGh<�h=Kub����       �8       K��R�}�(hKhiMhjh))��}�(h,h/h0M��h2h3h4hph<�h=Kub������       Z                     @>AU`�z�?�           8�@                                   �?�Ƀ aA�?�            pr@                                   �?0�!F��?W            �`@        ������������������������       �                    �@@                                   :@P���Q�??             Y@                                   L@�����?             E@                                 @4@��p\�?            �D@                                  �? ��WV�?             :@       	       
                   �B@P���Q�?             4@       ������������������������       �                     .@                                  �,@z�G�z�?             @                                  D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                    �?�r����?	             .@        ������������������������       �                      @                                   6@8�Z$���?             *@        ������������������������       �                     �?                                   �?�8��8��?             (@                                 �E@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                   @ _�@�Y�?"             M@        ������������������������       �                     �?        ������������������������       �        !            �L@               Q                     �?������?k            @d@              N                   �J@X�Cc�?>            �X@               !                   �9@��Zy�?/            �S@        ������������������������       �                     @        "       K                    �?)O���?*             R@       #       F                 ���X@��:c���?'            �P@       $       ?                   �G@��B����?              J@       %       *                    <@���Q��?             D@        &       )                    �?z�G�z�?             $@       '       (                   �6@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        +       0                    �?������?             >@        ,       /                    �?؇���X�?             @       -       .                   �A@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        1       6                 `f�;@8����?             7@        2       3                 03k:@      �?             @        ������������������������       �                     �?        4       5                 �|�?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        7       >                    D@���y4F�?             3@        8       9                 �|Y=@���Q��?             $@        ������������������������       �                      @        :       ;                 0�?D@      �?              @        ������������������������       �                      @        <       =                   @K@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        @       E                 �5L@�8��8��?             (@       A       D                   �I@r�q��?             @       B       C                 �̜D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        G       J                    �?z�G�z�?             .@       H       I                 p�w@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        L       M                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        O       P                   �R@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        R       S                    %@     ��?-             P@        ������������������������       �                     @        T       Y                    4@ _�@�Y�?(             M@        U       V                   �2@      �?             @        ������������������������       �                      @        W       X                   �'@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        $             K@        [       �                    �?�3�E���?            z@        \       q                    �?��S���?J             ^@        ]       p                 X�,A@     ��?             H@       ^       c                    (@�r����?            �F@        _       b                 `�@1@���Q��?             @        `       a                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        d       m                    �?ףp=
�?             D@        e       f                 �|Y=@r�q��?             (@        ������������������������       �                     @        g       l                    �?�q�q�?             @       h       k                    �?z�G�z�?             @       i       j                 ��%@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        n       o                 ���@@4և���?             <@        ������������������������       �                      @        ������������������������       �                     :@        ������������������������       �                     @        r       �                    �?<ݚ�?-             R@       s       |                   �:@�n_Y�K�?            �C@        t       u                 ��y@�	j*D�?
             *@        ������������������������       �                     �?        v       y                   �6@      �?	             (@       w       x                 ؼC1@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        z       {                 �0@      �?             @       ������������������������       �                      @        ������������������������       �                      @        }       �                 03�-@�θ�?             :@       ~                        ���@؇���X�?             5@        ������������������������       �                      @        �       �                   @@�θ�?             *@        �       �                 �|=@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        �       �                 �|Y=@�����H�?             "@        �       �                    <@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�FVQ&�?            �@@       �       �                   `3@�>����?             ;@       �       �                 ��(@ ��WV�?             :@       �       �                 X��A@�X�<ݺ?             2@       �       �                 ���@��S�ۿ?	             .@        ������������������������       �                     @        ������������������������       ������H�?             "@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?��A��?�            �r@        �       �                    �?����X�?             @        ������������������������       �                     @        �       �                 ��!>@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                 pff/@x{&�cn�?�            r@       �       �                    �?��?��:�?�            �j@        �       �                 ���@*;L]n�?             >@        ������������������������       �                     @        �       �                   �3@��+7��?             7@        ������������������������       �                     @        �       �                 �|�=@�KM�]�?             3@       ������������������������       �        
             ,@        �       �                   &@���Q��?             @        ������������������������       �                      @        �       �                   @C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �?�@85�}C�?r            �f@       �       �                   �@X;��?:            @V@       �       �                    7@����˵�?(            �M@        ������������������������       �                     6@        �       �                   �8@�L���?            �B@        �       �                 `fF@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @@@ >�֕�?            �A@        �       �                   �?@�t����?             1@       �       �                 pf�@      �?             0@       ������������������������       �                     "@        �       �                 �|�<@؇���X�?             @        ������������������������       �                      @        �       �                 �|Y>@z�G�z�?             @       ������������������������       �      �?             @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     >@        �       �                   �;@��E�B��?8            �W@        �       �                   �:@4�2%ޑ�?            �A@       �       �                 0S5 @     ��?             @@       �       �                 @3�@�E��ӭ�?             2@        �       �                   �4@؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        �       �                   �4@���|���?             &@       �       �                    1@և���X�?             @        ������������������������       �                      @        �       �                   �2@z�G�z�?             @        ������������������������       �                     @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        
             ,@        ������������������������       �                     @        �       �                 @3�@ ,��-�?"            �M@        �       �                   �?@      �?              @        �       �                   �=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    ?@`'�J�?            �I@       �       �                 ��) @      �?             @@        ������������������������       �        	             ,@        �       �                 pf� @�����H�?	             2@        ������������������������       �                     �?        �       �                 �|�=@�IєX�?             1@       ������������������������       �                     0@        ������������������������       �                     �?        ������������������������       �                     3@        �       �                   �6@      �?1             S@        �       �                    �? 	��p�?             =@       �       �                    0@�KM�]�?
             3@        ������������������������       �                     �?        �       �                    �?�X�<ݺ?	             2@       �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �                 @3�2@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �        	             $@        �       �                    �?Z�K�D��?            �G@        �       �                   @@@r�q��?             8@       �       �                 ��1@�G�z��?             4@        �       �                 �|�;@      �?              @        ������������������������       �                     �?        �       �                 @3�/@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 �T)D@�q�q�?             (@        ������������������������       �                     @        �       �                    ;@և���X�?             @        ������������������������       �                      @        �       �                 �|�>@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �̜2@�㙢�c�?             7@        �       �                    A@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �                           @�}�+r��?             3@       ������������������������       �                     1@                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �*       h�h))��}�(h,h/h0MKK��h2h3h4hVh<�h=Kub������������.���|�?ӣ���?'u_�?~ylE�p�?�3�τ?�?�����?              �?�������?ffffff�?�a�a�?=��<���?��+Q��?�]�ڕ��?;�;��?O��N���?�������?ffffff�?              �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�?�������?              �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?      �?                      �?      �?        �{a���?#,�4�r�?      �?                      �?B{	�%��?{	�%���?%I�$I��?�m۶m��?� � �?\��[���?      �?        9��8���?��8��8�?*g���?�1���?O��N���?ى�؉��?333333�?�������?�������?�������?�q�q�?9��8���?      �?                      �?              �?wwwwww�?�?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?                      �?      �?        d!Y�B�?8��Moz�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?6��P^C�?(������?333333�?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?�������?      �?      �?      �?                      �?      �?        �������?�������?      �?                      �?ffffff�?�������?      �?                      �?     ��?      �?              �?#,�4�r�?�{a���?      �?      �?      �?              �?      �?              �?      �?              �?        ;�;��?ى�؉��?�?�������?      �?      �?�?�������?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?      �?        �$I�$I�?n۶m۶�?      �?                      �?      �?        �q�q�?��8��8�?;�;��?ى�؉��?;�;��?vb'vb'�?      �?              �?      �?      �?      �?              �?      �?              �?      �?      �?                      �?ى�؉��?�؉�؉�?۶m۶m�?�$I�$I�?      �?        ى�؉��?�؉�؉�?      �?      �?      �?        UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?      �?      �?                      �?      �?        �������?333333�?      �?                      �?>����?|���?�Kh/��?h/�����?O��N���?;�;��?��8��8�?�q�q�?�������?�?      �?        �q�q�?�q�q�?      �?              �?                      �?      �?        ��g�`�?�g�`�|�?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?        �������?���I��?����?��χ��?""""""�?�������?              �?zӛ����?Y�B��?              �?�k(���?(�����?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �}�K�`�?������?�u�{���?�E(B�?W'u_�?��/���?      �?        }���g�?L�Ϻ��?      �?      �?              �?      �?        ��+��+�?�A�A�?<<<<<<�?�?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?      �?      �?      �?                      �?      �?              �?        �l�w6��?AL� &W�?�������?�A�A�?      �?      �?�q�q�?r�q��?۶m۶m�?�$I�$I�?      �?      �?      �?        ]t�E]�?F]t�E�?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?      �?      �?              �?                      �?[4���?'u_[�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�?      �?      �?      �?        �q�q�?�q�q�?              �?�?�?      �?                      �?      �?              �?      �?������?�{a���?�k(���?(�����?              �?��8��8�?�q�q�?�q�q�?�q�q�?      �?        �������?�������?              �?      �?              �?              �?        R�٨�l�?]AL� &�?UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?              �?333333�?�������?      �?                      �?              �?�7��Mo�?d!Y�B�?      �?      �?              �?      �?        �5��P�?(�����?      �?              �?      �?              �?      �?        �       ubhhubehhub.